CircuitMaker Text
5.6
Probes: 1
U2_6
Transient Analysis
0 353 192 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 130 10
176 79 1918 540
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
22
11 Signal Gen~
195 33 240 0 64 64
0 6 7 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1073741824 1073741824
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 2 2 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/4V
-15 -30 13 -22
2 V3
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(2 2 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5130 0 0
2
5.89861e-315 5.39306e-315
0
8 Op-Amp5~
219 299 87 0 5 11
0 18 17 19 2 16
0
0 0 848 0
5 AD820
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
391 0 0
2
5.89861e-315 5.38788e-315
0
11 Signal Gen~
195 33 86 0 64 64
0 13 7 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1127481344 1127481344
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 180 180 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
6 0/360V
-21 -30 21 -22
2 V2
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(180 180 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3124 0 0
2
5.89861e-315 5.37752e-315
0
7 Ground~
168 248 158 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3421 0 0
2
5.89861e-315 5.36716e-315
0
2 +V
167 299 58 0 1 3
0 19
0
0 0 53616 0
4 3.3v
-13 -13 15 -5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8157 0 0
2
5.89861e-315 5.3568e-315
0
7 Ground~
168 299 110 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5572 0 0
2
5.89861e-315 5.34643e-315
0
7 Ground~
168 300 264 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8901 0 0
2
5.89861e-315 5.32571e-315
0
2 +V
167 300 212 0 1 3
0 12
0
0 0 53616 0
4 3.3v
-13 -13 15 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7361 0 0
2
5.89861e-315 5.30499e-315
0
7 Ground~
168 249 312 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4747 0 0
2
5.89861e-315 5.26354e-315
0
8 Op-Amp5~
219 300 241 0 5 11
0 3 4 12 2 11
0
0 0 848 0
5 AD820
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
972 0 0
2
5.89861e-315 0
0
11 Resistor:A~
219 300 31 0 2 5
0 17 16
0
0 0 880 0
2 3k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3472 0 0
2
5.89861e-315 5.44228e-315
0
11 Resistor:A~
219 248 127 0 3 5
0 2 18 -1
0
0 0 880 90
2 3k
9 -1 23 7
2 R3
9 -12 23 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9998 0 0
2
5.89861e-315 5.43969e-315
0
11 Resistor:A~
219 219 93 0 2 5
0 14 18
0
0 0 880 0
4 124k
-16 17 12 25
2 R2
-10 7 4 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3536 0 0
2
5.89861e-315 5.4371e-315
0
11 Resistor:A~
219 219 81 0 2 5
0 15 17
0
0 0 880 0
4 124k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4597 0 0
2
5.89861e-315 5.43451e-315
0
11 Resistor:A~
219 149 81 0 2 5
0 7 15
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3835 0 0
2
5.89861e-315 5.43192e-315
0
11 Resistor:A~
219 149 93 0 2 5
0 13 14
0
0 0 880 0
4 224k
-16 17 12 25
2 R7
-10 7 4 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3670 0 0
2
5.89861e-315 5.42933e-315
0
11 Resistor:A~
219 249 281 0 3 5
0 2 3 -1
0
0 0 880 90
4 270k
9 -1 37 7
3 R12
6 -12 27 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5616 0 0
2
5.89861e-315 5.42414e-315
0
11 Resistor:A~
219 301 185 0 2 5
0 4 11
0
0 0 880 0
4 270k
-14 -14 14 -6
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9323 0 0
2
5.89861e-315 5.41896e-315
0
11 Resistor:A~
219 149 247 0 2 5
0 6 8
0
0 0 880 0
4 224k
-16 17 12 25
2 R5
-10 7 4 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
317 0 0
2
5.89861e-315 5.41378e-315
0
11 Resistor:A~
219 149 235 0 2 5
0 7 9
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3108 0 0
2
5.89861e-315 5.4086e-315
0
11 Resistor:A~
219 219 235 0 2 5
0 9 4
0
0 0 880 0
4 124k
-14 -14 14 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4299 0 0
2
5.89861e-315 5.40342e-315
0
11 Resistor:A~
219 219 247 0 2 5
0 8 3
0
0 0 880 0
4 124k
-15 18 13 26
3 R10
-13 7 8 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9672 0 0
2
5.89861e-315 5.39824e-315
0
27
2 0 3 0 0 4096 0 22 0 0 13 2
237 247
249 247
2 0 4 0 0 4096 0 21 0 0 14 2
237 235
249 235
0 0 5 0 0 0 0 0 0 0 0 2
153 224
153 224
1 1 6 0 0 12416 0 1 19 0 0 6
64 235
85 235
85 255
109 255
109 247
131 247
2 1 7 0 0 12288 0 1 20 0 0 4
64 245
92 245
92 235
131 235
2 1 8 0 0 4224 0 19 22 0 0 2
167 247
201 247
1 2 9 0 0 4224 0 21 20 0 0 2
201 235
167 235
0 0 10 0 0 0 0 0 0 0 0 2
153 70
153 70
0 0 7 0 0 4224 0 0 0 17 5 2
69 91
69 245
2 5 11 0 0 8320 0 18 10 0 0 4
319 185
353 185
353 241
318 241
1 3 12 0 0 4224 0 8 10 0 0 2
300 221
300 228
1 4 2 0 0 4096 0 7 10 0 0 2
300 258
300 254
2 1 3 0 0 8320 0 17 10 0 0 3
249 263
249 247
282 247
1 2 4 0 0 8320 0 18 10 0 0 4
283 185
249 185
249 235
282 235
1 1 2 0 0 4224 0 9 17 0 0 2
249 306
249 299
1 1 13 0 0 12416 0 3 16 0 0 6
64 81
85 81
85 101
109 101
109 93
131 93
2 1 7 0 0 0 0 3 15 0 0 4
64 91
92 91
92 81
131 81
2 1 14 0 0 4224 0 16 13 0 0 2
167 93
201 93
1 2 15 0 0 4224 0 14 15 0 0 2
201 81
167 81
2 5 16 0 0 8320 0 11 2 0 0 4
318 31
352 31
352 87
317 87
0 1 17 0 0 4224 0 0 11 26 0 3
248 81
248 31
282 31
2 0 18 0 0 4096 0 12 0 0 25 2
248 109
248 93
1 3 19 0 0 4224 0 5 2 0 0 2
299 67
299 74
1 4 2 0 0 0 0 6 2 0 0 2
299 104
299 100
1 2 18 0 0 4224 0 2 13 0 0 2
281 93
237 93
2 2 17 0 0 0 0 2 14 0 0 2
281 81
237 81
1 1 2 0 0 0 0 4 12 0 0 2
248 152
248 145
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.1 0.0004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
