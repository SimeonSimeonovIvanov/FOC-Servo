CircuitMaker Text
5.6
Probes: 1
U3_1
Transient Analysis
0 671 91 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 79 1918 469
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.576596 0.500000
344 175 2086 716
9961490 0
0
6 Title:
5 Name:
0
0
0
24
8 Op-Amp5~
219 621 98 0 5 11
0 3 4 9 2 8
0
0 0 848 0
7 MAX4212
10 10 59 18
2 U3
12 -12 26 -4
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
7 SOT23-5
11

0 3 4 5 2 1 3 4 5 2
1 0
88 0 0 256 1 0 0 0
1 U
6369 0 0
2
43307 4
0
2 +V
167 492 147 0 1 3
0 5
0
0 0 53616 90
5 1.65V
-40 -6 -5 2
3 V11
-46 -15 -25 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9172 0 0
2
43307 3
0
11 Signal Gen~
195 421 96 0 64 64
0 7 6 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1092616192
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 1000 0 10 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -10/10V
-25 -30 24 -22
3 V12
-10 -40 11 -32
0
0
37 %D %1 %2 DC 0 SIN(0 10 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
43307 2
0
7 Ground~
168 621 132 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
43307 1
0
2 +V
167 621 63 0 1 3
0 9
0
0 0 53616 0
3 10V
-10 -16 11 -8
3 V13
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7678 0 0
2
43307 0
0
7 Ground~
168 69 156 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
961 0 0
2
43307 0
0
11 Signal Gen~
195 30 103 0 64 64
0 11 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1092616192
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 70
20
1 1000 0 10 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -10/10V
-25 -30 24 -22
2 V4
-8 -40 6 -32
0
0
37 %D %1 %2 DC 0 SIN(0 10 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3178 0 0
2
43307 1
0
7 Ground~
168 129 156 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3409 0 0
2
43307 2
0
2 +V
167 206 141 0 1 3
0 12
0
0 0 54128 90
5 3.30V
-39 -5 -4 3
2 V3
-29 -15 -15 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3951 0 0
2
43307 3
0
2 +V
167 210 88 0 1 3
0 14
0
0 0 54128 90
5 1.65V
-38 -6 -3 2
2 V2
-28 -16 -14 -8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8885 0 0
2
43307 4
0
7 Ground~
168 303 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3780 0 0
2
43307 5
0
2 +V
167 303 64 0 1 3
0 15
0
0 0 54128 0
4 3.3V
-12 -16 16 -8
2 V1
-5 -26 9 -18
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9265 0 0
2
43307 6
0
8 Op-Amp5~
219 303 92 0 5 11
0 13 17 15 2 16
0
0 0 848 0
10 LM6132A/NS
8 6 78 14
3 U1B
9 -14 30 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
9442 0 0
2
43307 7
0
11 Resistor:A~
219 552 145 0 3 5
0 5 3 1
0
0 0 880 0
2 1k
-6 21 8 29
3 R10
-9 8 12 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9424 0 0
2
43307 9
0
11 Resistor:A~
219 494 98 0 2 5
0 6 7
0
0 0 880 90
3 10k
5 0 26 8
3 R11
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9968 0 0
2
43307 8
0
11 Resistor:A~
219 584 68 0 2 5
0 4 8
0
0 0 880 90
2 1k
8 0 22 8
3 R12
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9281 0 0
2
43307 7
0
11 Resistor:A~
219 553 92 0 2 5
0 7 4
0
0 0 880 0
5 7.40k
-17 -14 18 -6
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8464 0 0
2
43307 6
0
11 Resistor:A~
219 553 104 0 2 5
0 6 3
0
0 0 880 0
5 7.40k
-17 16 18 24
3 R14
-10 6 11 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
43307 5
0
11 Resistor:A~
219 103 98 0 2 5
0 11 10
0
0 0 880 0
4 6.2k
-12 8 16 16
2 R6
-11 -14 3 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3171 0 0
2
43307 8
0
11 Resistor:A~
219 129 124 0 3 5
0 2 10 -1
0
0 0 880 90
4 1.1k
8 0 36 8
2 R5
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4139 0 0
2
43307 9
0
11 Resistor:A~
219 246 139 0 3 5
0 12 13 1
0
0 0 880 0
3 51k
-14 20 7 28
2 R4
-11 10 3 18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6435 0 0
2
43307 10
0
11 Resistor:A~
219 247 98 0 2 5
0 10 13
0
0 0 880 0
3 51k
-14 20 7 28
2 R3
-11 10 3 18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5283 0 0
2
43307 11
0
11 Resistor:A~
219 303 29 0 2 5
0 17 16
0
0 0 880 0
3 51k
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6874 0 0
2
43307 12
0
11 Resistor:A~
219 247 86 0 3 5
0 14 17 1
0
0 0 880 0
3 51k
-15 -15 6 -7
2 R1
-12 -25 2 -17
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5305 0 0
2
43307 13
0
26
2 0 3 0 0 8336 0 14 0 0 3 3
570 145
584 145
584 104
1 0 4 0 0 4112 0 16 0 0 10 2
584 86
584 92
2 1 3 0 0 16 0 18 1 0 0 2
571 104
603 104
1 1 5 0 0 4240 0 2 14 0 0 2
503 145
534 145
2 0 6 0 0 4112 0 3 0 0 7 4
452 101
475 101
475 124
494 124
1 0 7 0 0 4112 0 3 0 0 8 4
452 91
475 91
475 69
493 69
1 1 6 0 0 12432 0 18 15 0 0 5
535 104
525 104
525 124
494 124
494 116
1 2 7 0 0 12432 0 17 15 0 0 7
535 92
525 92
525 69
493 69
493 69
494 69
494 80
2 5 8 0 0 8336 0 16 1 0 0 5
584 50
584 38
672 38
672 98
639 98
2 2 4 0 0 4240 0 17 1 0 0 2
571 92
603 92
1 4 2 0 0 4112 0 4 1 0 0 2
621 126
621 111
3 1 9 0 0 4240 0 1 5 0 0 2
621 85
621 72
1 0 10 0 0 4224 0 22 0 0 17 2
229 98
129 98
1 1 11 0 0 4224 0 7 19 0 0 2
61 98
85 98
1 2 2 0 0 4224 0 6 7 0 0 3
69 150
69 108
61 108
1 1 2 0 0 0 0 8 20 0 0 2
129 150
129 142
2 2 10 0 0 0 0 20 19 0 0 3
129 106
129 98
121 98
1 1 12 0 0 4224 0 9 21 0 0 2
217 139
228 139
2 0 13 0 0 4096 0 22 0 0 20 2
265 98
273 98
2 1 13 0 0 8320 0 21 13 0 0 4
264 139
273 139
273 98
285 98
1 1 14 0 0 4224 0 10 24 0 0 2
221 86
229 86
1 3 15 0 0 4224 0 12 13 0 0 2
303 73
303 79
1 4 2 0 0 0 0 11 13 0 0 2
303 112
303 105
2 5 16 0 0 8320 0 23 13 0 0 4
321 29
354 29
354 92
321 92
1 0 17 0 0 8320 0 23 0 0 26 3
285 29
273 29
273 86
2 2 17 0 0 0 0 24 13 0 0 2
265 86
285 86
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
