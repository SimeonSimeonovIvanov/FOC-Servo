CircuitMaker Text
5.6
Probes: 4
U1A_1
AC Analysis
0 279 93 65280
U1A_1
DC Sweep
0 279 93 65280
U1A_1
Fourier Analysis
0 279 93 65280
U1A_1
Transient Analysis
0 307 113 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 230 10
176 79 1918 1019
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 2 1
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
13
10 Capacitor~
219 274 46 0 2 5
0 4 3
0
0 0 848 0
4 22pF
-13 -18 15 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
5551 0 0
2
42785.8 0
0
2 +V
167 155 135 0 1 3
0 5
0
0 0 53616 90
5 1.55V
-23 -16 12 -8
2 V1
-6 -28 8 -20
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6986 0 0
2
42785.8 7
0
7 Ground~
168 99 173 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8745 0 0
2
42785.8 6
0
11 Signal Gen~
195 58 150 0 64 64
0 6 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1182938454 0 1065353216
0 897988541 897988541 939239554 947628162 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 16666.7 0 1 0 1e-06 1e-06 3e-05 6e-05 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/1V
-13 -30 15 -22
2 V3
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 PULSE(0 1 0 1u 1u 30u 60u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9592 0 0
2
42785.8 5
0
7 Ground~
168 246 165 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8748 0 0
2
42785.8 4
0
8 Op-Amp5~
219 246 139 0 5 11
0 8 4 9 2 3
0
0 0 848 0
6 OP284E
12 -25 54 -17
3 U1A
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
7168 0 0
2
42785.8 3
0
2 +V
167 246 112 0 1 3
0 9
0
0 0 53616 0
4 3.3V
-13 -14 15 -6
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
631 0 0
2
42785.8 2
0
2 +V
167 130 77 0 1 3
0 7
0
0 0 53616 0
4 3.3V
-13 -14 15 -6
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9466 0 0
2
42785.8 1
0
5 SAVE-
218 305 137 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3266 0 0
2
42785.8 0
0
11 Resistor:A~
219 217 186 0 2 5
0 6 8
0
0 0 880 90
4 3.3k
-32 1 -4 9
2 R2
-28 -10 -14 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7693 0 0
2
42785.8 11
0
11 Resistor:A~
219 245 76 0 2 5
0 4 3
0
0 0 880 0
4 3.3k
-13 -14 15 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3723 0 0
2
42785.8 10
0
11 Resistor:A~
219 185 133 0 3 5
0 5 4 1
0
0 0 880 0
4 3.3k
-13 -14 15 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3440 0 0
2
42785.8 9
0
11 Resistor:A~
219 185 145 0 3 5
0 7 8 1
0
0 0 880 0
4 3.3k
-15 14 13 22
2 R3
-12 5 2 13
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6263 0 0
2
42785.8 8
0
14
2 0 3 0 0 8192 0 1 0 0 8 3
283 46
305 46
305 76
1 0 4 0 0 4112 0 1 0 0 9 3
265 46
217 46
217 76
1 1 5 0 0 4224 0 2 12 0 0 2
166 133
167 133
1 1 6 0 0 12416 0 4 10 0 0 5
89 145
119 145
119 225
217 225
217 204
1 1 7 0 0 8320 0 13 8 0 0 3
167 145
130 145
130 86
2 1 2 0 0 8320 0 4 3 0 0 3
89 155
99 155
99 167
2 0 8 0 0 4096 0 10 0 0 11 2
217 168
217 145
2 5 3 0 0 8320 0 11 6 0 0 4
263 76
305 76
305 139
264 139
1 0 4 0 0 8320 0 11 0 0 10 3
227 76
217 76
217 133
2 2 4 0 0 0 0 12 6 0 0 2
203 133
228 133
2 1 8 0 0 4224 0 13 6 0 0 2
203 145
228 145
1 4 2 0 0 0 0 5 6 0 0 2
246 159
246 152
1 3 9 0 0 4224 0 7 6 0 0 2
246 121
246 126
0 0 10 0 0 0 0 0 0 0 0 2
30 94
30 94
0
0
2065 2 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.003 1.2e-06 1.2e-06
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
