CircuitMaker Text
5.6
Probes: 1
C1_2
Transient Analysis
0 472 120 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 79 1918 540
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
28
2 +V
167 220 166 0 1 3
0 17
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V1
-7 -10 7 -2
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9604 0 0
2
43307 0
0
7 Ground~
168 178 187 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7518 0 0
2
43307 0
0
2 +V
167 220 89 0 1 3
0 18
0
0 0 53616 0
3 15V
-10 -16 11 -8
3 V13
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4832 0 0
2
43307 27
0
8 Op-Amp5~
219 220 124 0 5 11
0 3 16 18 17 8
0
0 0 848 0
7 MAX4212
10 10 59 18
2 U3
12 -12 26 -4
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
7 SOT23-5
11

0 3 4 5 2 1 3 4 5 2
1 0
88 0 0 256 1 0 0 0
1 U
6798 0 0
2
43307 24
0
11 Signal Gen~
195 31 122 0 64 64
0 4 5 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1073741824 1070805811 1068289229
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 2 1.65 1.35 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 300m/3V
-25 -30 24 -22
2 V7
-8 -40 6 -32
0
0
41 %D %1 %2 DC 0 SIN(1.65 1.35 2 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3336 0 0
2
43307 23
0
2 +V
167 423 153 0 1 3
0 12
0
0 0 53616 180
4 -15V
-14 0 14 8
2 V9
-7 -10 7 -2
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8370 0 0
2
43307 22
0
2 +V
167 423 102 0 1 3
0 13
0
0 0 53616 0
4 +15V
-12 -14 16 -6
2 V8
-5 -24 9 -16
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3910 0 0
2
43307 21
0
7 Ground~
168 319 184 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
316 0 0
2
43307 20
0
2 +V
167 364 276 0 1 3
0 10
0
0 0 53616 180
4 -15V
-13 1 15 9
2 V6
-6 -9 8 -1
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
536 0 0
2
43307 19
0
7 N-JFET~
219 386 176 0 3 7
0 11 9 2
0
0 0 848 0
6 2N4393
12 0 54 8
2 Q1
26 -10 40 -2
0
0
14 %D %1 %2 %3 %M
0
0
5 TO-18
7

0 2 3 1 2 3 1 0
74 0 0 0 1 0 0 0
1 Q
4460 0 0
2
43307 18
0
7 Ground~
168 394 272 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3260 0 0
2
43307 17
0
8 Op-Amp5~
219 423 124 0 5 11
0 11 7 13 12 6
0
0 0 848 0
5 TL082
9 -12 44 -4
3 U4A
16 -22 37 -14
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 2 0
1 U
5156 0 0
2
43307 16
0
7 Ground~
168 339 272 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3133 0 0
2
43307 15
0
14 Opto Isolator~
173 305 239 0 4 9
0 15 2 9 2
0
0 0 880 0
6 OP4N25
-20 20 22 28
2 U2
-6 -29 8 -21
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 0
88 0 0 0 1 0 0 0
1 U
5523 0 0
2
43307 14
0
11 Signal Gen~
195 31 232 0 64 64
0 14 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1056964608 0 1079194419
0 814313567 814313567 1065353216 1073741824 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 258
20
0 0.5 0 3.3 0 1e-09 1e-09 1 2 0
0 0 0 0 0 0 0 0 0 0
0
0 0 1360 0
6 0/3.3V
-21 -30 21 -22
2 V5
-8 -40 6 -32
4 F/!B
-13 -44 15 -36
0
38 %D %1 %2 DC 0 PULSE(0 3.3 0 1n 1n 1 2)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3746 0 0
2
43307 13
0
7 Ground~
168 262 270 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5668 0 0
2
43307 12
0
10 Capacitor~
219 423 34 0 2 5
0 7 6
0
0 0 848 0
6 0.01uF
-21 -18 21 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
5368 0 0
2
43307 0
0
11 Resistor:A~
219 152 130 0 2 5
0 4 3
0
0 0 880 0
3 10k
-10 16 11 24
3 R14
-10 6 11 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8293 0 0
2
43307 11
0
11 Resistor:A~
219 152 118 0 2 5
0 5 16
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3232 0 0
2
43307 10
0
11 Resistor:A~
219 178 91 0 2 5
0 16 8
0
0 0 880 90
3 33k
5 0 26 8
3 R12
9 -10 30 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6644 0 0
2
43307 9
0
11 Resistor:A~
219 93 124 0 2 5
0 4 5
0
0 0 880 90
3 10k
5 0 26 8
3 R11
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4978 0 0
2
43307 8
0
11 Resistor:A~
219 178 155 0 3 5
0 2 3 -1
0
0 0 880 90
3 33k
7 0 28 8
3 R10
7 -10 28 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9207 0 0
2
43307 7
0
11 Resistor:A~
219 423 63 0 2 5
0 7 6
0
0 0 880 0
3 10k
-12 9 9 17
3 R17
-14 -14 7 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6998 0 0
2
43307 6
0
11 Resistor:A~
219 366 118 0 2 5
0 8 7
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R16
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3175 0 0
2
43307 5
0
11 Resistor:A~
219 366 130 0 2 5
0 8 11
0
0 0 880 0
3 10k
-11 18 10 26
3 R15
-11 8 10 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3378 0 0
2
43307 4
0
11 Resistor:A~
219 319 154 0 3 5
0 2 8 -1
0
0 0 880 90
3 10k
-28 1 -7 9
2 R9
-25 -9 -11 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
922 0 0
2
43307 3
0
11 Resistor:A~
219 364 201 0 3 5
0 10 9 1
0
0 0 880 90
3 20k
7 0 28 8
2 R8
10 -10 24 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6891 0 0
2
43307 2
0
11 Resistor:A~
219 254 227 0 2 5
0 15 14
0
0 0 880 180
3 100
-11 -14 10 -6
2 R7
-8 -24 6 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5407 0 0
2
43307 1
0
34
1 1 2 0 0 4096 0 2 22 0 0 2
178 181
178 173
2 0 3 0 0 4096 0 22 0 0 28 2
178 137
178 130
0 1 4 0 0 8320 0 0 5 29 0 4
93 150
69 150
69 117
62 117
2 0 5 0 0 8320 0 5 0 0 30 4
62 127
80 127
80 95
92 95
2 0 6 0 0 4096 0 17 0 0 15 3
432 34
471 34
471 63
1 0 7 0 0 8192 0 17 0 0 16 3
414 34
395 34
395 63
0 0 8 0 0 8192 0 0 0 31 8 3
271 123
271 124
319 124
2 0 8 0 0 0 0 26 0 0 20 3
319 136
319 124
340 124
1 0 2 0 0 4096 0 16 0 0 24 2
262 264
262 251
3 0 9 0 0 8320 0 14 0 0 12 4
331 227
338 227
338 176
364 176
1 1 10 0 0 4224 0 9 27 0 0 2
364 261
364 219
2 2 9 0 0 0 0 27 10 0 0 3
364 183
364 176
373 176
1 3 2 0 0 4096 0 11 10 0 0 2
394 266
394 194
0 1 11 0 0 4224 0 0 10 22 0 2
394 130
394 158
2 5 6 0 0 8320 0 23 12 0 0 4
441 63
471 63
471 124
441 124
1 0 7 0 0 8320 0 23 0 0 21 3
405 63
394 63
394 118
4 1 12 0 0 4224 0 12 6 0 0 2
423 137
423 138
3 1 13 0 0 0 0 12 7 0 0 2
423 111
423 111
1 1 2 0 0 0 0 8 26 0 0 2
319 178
319 172
1 1 8 0 0 0 0 25 24 0 0 4
348 130
340 130
340 118
348 118
2 2 7 0 0 0 0 24 12 0 0 2
384 118
405 118
2 1 11 0 0 0 0 25 12 0 0 2
384 130
405 130
1 4 2 0 0 0 0 13 14 0 0 3
339 266
339 251
331 251
2 2 2 0 0 4224 0 14 15 0 0 4
277 251
85 251
85 237
62 237
1 2 14 0 0 4224 0 15 28 0 0 2
62 227
236 227
1 1 15 0 0 4224 0 28 14 0 0 2
272 227
277 227
1 0 16 0 0 4096 0 20 0 0 32 2
178 109
178 118
2 1 3 0 0 4224 0 18 4 0 0 2
170 130
202 130
1 1 4 0 0 128 0 18 21 0 0 5
134 130
124 130
124 150
93 150
93 142
1 2 5 0 0 128 0 19 21 0 0 7
134 118
124 118
124 95
92 95
92 95
93 95
93 106
2 5 8 0 0 8320 0 20 4 0 0 5
178 73
178 64
271 64
271 124
238 124
2 2 16 0 0 4224 0 19 4 0 0 2
170 118
202 118
1 4 17 0 0 4224 0 1 4 0 0 2
220 151
220 137
3 1 18 0 0 4224 0 4 3 0 0 2
220 111
220 98
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 4 0.002 0.002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
