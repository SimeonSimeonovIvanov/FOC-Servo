CircuitMaker Text
5.6
Probes: 2
C4_2
Operating Point
0 760 120 65280
C4_2
Transient Analysis
0 759 175 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 160 10
241 79 1918 470
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 0 1
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.575532 0.500000
409 175 2086 715
9961474 0
0
2 

2 

0
0
0
24
10 Op-Amp5:A~
219 266 83 0 5 11
0 13 11 14 2 12
0
0 0 848 0
5 AD820
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 0 0 0 0
1 U
6169 0 0
2
43356 0
0
10 Op-Amp5:A~
219 690 83 0 5 11
0 7 5 8 2 6
0
0 0 848 0
5 AD820
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 0 0 0 0
1 U
3362 0 0
2
43356 0
0
11 Signal Gen~
195 28 82 0 64 64
0 10 3 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1127481344 1127481344
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 180 180 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
6 0/360V
-21 -30 21 -22
2 V1
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(180 180 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4391 0 0
2
43356 15
0
7 Ground~
168 266 112 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8214 0 0
2
43356 13
0
2 +V
167 266 55 0 1 3
0 14
0
0 0 54128 0
2 5V
-6 -13 8 -5
2 V2
-6 -23 8 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7266 0 0
2
43356 12
0
10 Capacitor~
219 270 200 0 2 5
0 11 12
0
0 0 848 0
4 10nF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3947 0 0
2
43356 11
0
10 Capacitor~
219 188 44 0 2 5
0 13 2
0
0 0 848 90
4 10nF
12 0 40 8
2 C2
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5715 0 0
2
43356 10
0
7 Ground~
168 143 9 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5703 0 0
2
43356 9
0
7 Ground~
168 188 9 0 1 3
0 2
0
0 0 53360 180
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3511 0 0
2
43356 8
0
11 Signal Gen~
195 453 82 0 64 64
0 4 3 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1084227584 1073741824 1073741824
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 5 2 2 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/4V
-15 -30 13 -22
2 V3
-8 -40 6 -32
0
0
35 %D %1 %2 DC 0 SIN(2 2 5 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
9901 0 0
2
43356 7
0
7 Ground~
168 612 9 0 1 3
0 2
0
0 0 53360 180
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9115 0 0
2
43356 6
0
7 Ground~
168 567 9 0 1 3
0 2
0
0 0 53360 180
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5545 0 0
2
43356 5
0
10 Capacitor~
219 612 44 0 2 5
0 7 2
0
0 0 848 90
3 1nF
15 0 36 8
2 C3
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9700 0 0
2
43356 4
0
10 Capacitor~
219 694 200 0 2 5
0 5 6
0
0 0 848 0
3 1nF
-11 -18 10 -10
2 C4
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3905 0 0
2
43356 3
0
2 +V
167 690 55 0 1 3
0 8
0
0 0 54128 0
4 3.3V
-13 -13 15 -5
2 V4
-6 -23 8 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
976 0 0
2
43356 2
0
7 Ground~
168 690 112 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3676 0 0
2
43356 1
0
11 Resistor:A~
219 108 89 0 2 5
0 3 11
0
0 0 880 0
4 336k
-16 17 12 25
2 R1
-9 7 5 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6137 0 0
2
43356 23
0
11 Resistor:A~
219 108 77 0 2 5
0 10 13
0
0 0 880 0
4 336k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3458 0 0
2
43356 22
0
11 Resistor:A~
219 269 155 0 2 5
0 11 12
0
0 0 880 0
2 3k
-7 -14 7 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8160 0 0
2
43356 21
0
11 Resistor:A~
219 143 44 0 4 5
0 13 2 0 -1
0
0 0 880 90
2 3k
6 -2 20 6
2 R4
6 -12 20 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8874 0 0
2
43356 20
0
11 Resistor:A~
219 567 44 0 4 5
0 7 2 0 -1
0
0 0 880 90
2 1k
8 -2 22 6
2 R5
9 -12 23 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3791 0 0
2
43356 19
0
11 Resistor:A~
219 693 155 0 2 5
0 5 6
0
0 0 880 0
2 1k
-8 -14 6 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9555 0 0
2
43356 18
0
11 Resistor:A~
219 532 77 0 2 5
0 4 7
0
0 0 880 0
4 336k
-14 -14 14 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3215 0 0
2
43356 17
0
11 Resistor:A~
219 532 89 0 2 5
0 3 5
0
0 0 880 0
4 168k
-16 17 12 25
2 R8
-9 7 5 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7300 0 0
2
43356 16
0
31
0 0 3 0 0 8320 0 0 0 17 2 4
74 89
74 221
494 221
494 89
2 1 3 0 0 128 0 10 24 0 0 3
484 87
484 89
514 89
1 1 4 0 0 4224 0 10 23 0 0 2
484 77
514 77
1 0 5 0 0 4096 0 14 0 0 7 3
685 200
613 200
613 155
2 0 6 0 0 4096 0 14 0 0 6 3
703 200
760 200
760 155
5 2 6 0 0 8320 0 2 22 0 0 4
708 83
760 83
760 155
711 155
1 0 5 0 0 0 0 22 0 0 14 3
675 155
613 155
613 89
1 0 7 0 0 4096 0 13 0 0 15 2
612 53
612 77
1 0 7 0 0 0 0 21 0 0 15 2
567 62
567 77
1 2 2 0 0 4224 0 11 13 0 0 2
612 17
612 35
1 2 2 0 0 0 0 12 21 0 0 2
567 17
567 26
1 3 8 0 0 4224 0 15 2 0 0 2
690 64
690 70
4 1 2 0 0 0 0 2 16 0 0 4
690 96
690 95
690 95
690 106
2 2 5 0 0 4224 0 24 2 0 0 2
550 89
672 89
2 1 7 0 0 4224 0 23 2 0 0 2
550 77
672 77
0 0 9 0 0 0 0 0 0 0 0 2
594 66
594 66
2 1 3 0 0 128 0 3 17 0 0 4
59 87
60 87
60 89
90 89
1 1 10 0 0 4224 0 3 18 0 0 2
59 77
90 77
1 0 11 0 0 4096 0 6 0 0 22 3
261 200
189 200
189 155
2 0 12 0 0 4096 0 6 0 0 21 3
279 200
336 200
336 155
5 2 12 0 0 8320 0 1 19 0 0 4
284 83
336 83
336 155
287 155
1 0 11 0 0 0 0 19 0 0 29 3
251 155
189 155
189 89
1 0 13 0 0 4096 0 7 0 0 30 2
188 53
188 77
1 0 13 0 0 0 0 20 0 0 30 2
143 62
143 77
1 2 2 0 0 0 0 9 7 0 0 2
188 17
188 35
1 2 2 0 0 0 0 8 20 0 0 2
143 17
143 26
1 3 14 0 0 4224 0 5 1 0 0 2
266 64
266 70
4 1 2 0 0 0 0 1 4 0 0 2
266 96
266 106
2 2 11 0 0 4224 0 17 1 0 0 2
126 89
248 89
2 1 13 0 0 4224 0 18 1 0 0 2
126 77
248 77
0 0 15 0 0 0 0 0 0 0 0 2
170 66
170 66
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.8 0.0002 0.0002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
