CircuitMaker Text
5.6
Probes: 1
C5_2
Transient Analysis
0 434 146 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 220 10
176 79 1918 540
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 175 2086 645
9961490 0
0
2 

2 

0
0
0
19
10 Capacitor~
219 116 163 0 2 5
0 2 10
0
0 0 848 90
4 22nF
12 0 40 8
2 C1
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
513 0 0
2
43051.2 13
0
10 Capacitor~
219 171 164 0 2 5
0 2 11
0
0 0 848 90
4 22nF
12 0 40 8
2 C2
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8190 0 0
2
43051.2 12
0
10 Capacitor~
219 230 165 0 2 5
0 2 3
0
0 0 848 90
4 22nF
12 0 40 8
2 C3
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5209 0 0
2
43051.2 11
0
7 Ground~
168 116 186 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7239 0 0
2
43051.2 10
0
7 Ground~
168 171 186 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9474 0 0
2
43051.2 9
0
7 Ground~
168 230 186 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3783 0 0
2
43051.2 8
0
11 Signal Gen~
195 34 144 0 64 64
0 9 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1176256512 0 1084227584
0 814313567 814313567 944879383 953267991 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 10000 0 5 0 1e-09 1e-09 5e-05 0.0001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/5V
-15 -30 13 -22
2 V1
-8 -40 6 -32
0
0
41 %D %1 %2 DC 0 PULSE(0 5 0 1n 1n 50u 100u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5422 0 0
2
43051.2 7
0
7 Ground~
168 72 186 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8527 0 0
2
43051.2 6
0
10 Capacitor~
219 267 139 0 2 5
0 3 5
0
0 0 848 0
4 47nF
-16 -18 12 -10
2 C4
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
761 0 0
2
43051.2 5
0
2 +V
167 393 112 0 1 3
0 8
0
0 0 54128 0
2 7V
-7 -13 7 -5
2 V2
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7323 0 0
2
43051.2 4
0
8 Op-Amp5~
219 393 145 0 5 11
0 4 7 8 2 6
0
0 0 848 0
7 TCA0372
5 -18 54 -10
3 U1A
19 -28 40 -20
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP16
16

0 9 10 1 13 16 9 10 1 13
16 8 7 1 4 2 0
88 0 0 256 2 1 3 0
1 U
8543 0 0
2
43051.2 3
0
10 Capacitor~
219 400 35 0 2 5
0 7 6
0
0 0 848 0
6 0.15nF
-22 -18 20 -10
2 C5
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4240 0 0
2
43051.2 2
0
2 +V
167 365 153 0 1 3
0 4
0
0 0 54128 90
5 2.55V
-41 2 -6 10
2 V3
-31 -8 -17 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7857 0 0
2
43051.2 1
0
7 Ground~
168 393 171 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7255 0 0
2
43051.2 0
0
11 Resistor:A~
219 144 139 0 2 5
0 10 11
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R2
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7736 0 0
2
43051.2 18
0
11 Resistor:A~
219 200 139 0 2 5
0 11 3
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R3
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5435 0 0
2
43051.2 17
0
11 Resistor:A~
219 92 139 0 2 5
0 9 10
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R1
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3446 0 0
2
43051.2 16
0
11 Resistor:A~
219 307 139 0 2 5
0 5 7
0
0 0 880 0
2 1k
-6 -14 8 -6
2 R4
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3914 0 0
2
43051.2 15
0
11 Resistor:A~
219 400 75 0 2 5
0 7 6
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3948 0 0
2
43051.2 14
0
20
1 0 3 0 0 4240 0 9 0 0 16 2
258 139
230 139
1 4 2 0 0 4112 0 14 11 0 0 2
393 165
393 158
1 1 4 0 0 4240 0 13 11 0 0 2
376 151
375 151
2 1 5 0 0 4240 0 9 18 0 0 2
276 139
289 139
2 0 6 0 0 4112 0 12 0 0 10 3
409 35
454 35
454 75
1 0 7 0 0 4112 0 12 0 0 7 3
391 35
346 35
346 75
1 0 7 0 0 8336 0 19 0 0 8 3
382 75
346 75
346 139
2 2 7 0 0 16 0 18 11 0 0 2
325 139
375 139
1 3 8 0 0 4240 0 10 11 0 0 2
393 121
393 132
5 2 6 0 0 8336 0 11 19 0 0 4
411 145
454 145
454 75
418 75
1 2 2 0 0 4240 0 8 7 0 0 3
72 180
72 149
65 149
1 1 9 0 0 4240 0 7 17 0 0 2
65 139
74 139
1 1 2 0 0 16 0 6 3 0 0 2
230 180
230 174
1 1 2 0 0 16 0 5 2 0 0 2
171 180
171 173
1 1 2 0 0 16 0 4 1 0 0 2
116 180
116 172
2 2 3 0 0 16 0 16 3 0 0 3
218 139
230 139
230 156
2 0 10 0 0 4112 0 1 0 0 20 2
116 154
116 139
2 0 11 0 0 4112 0 2 0 0 19 2
171 155
171 139
2 1 11 0 0 4240 0 15 16 0 0 2
162 139
182 139
2 1 10 0 0 4240 0 17 15 0 0 2
110 139
126 139
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.002 2e-06 2e-06
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
