CircuitMaker Text
5.6
Probes: 1
R2_2
Transient Analysis
0 221 93 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
528 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 2 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
696 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
8
8 Op-Amp5~
219 176 92 0 5 11
0 5 7 3 2 6
0
0 0 848 0
10 LM6132A/NS
8 6 78 14
3 U1A
9 -14 30 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 83045552
88 0 0 256 2 1 1 0
1 U
4747 0 0
2
43302.6 0
0
2 +V
167 176 64 0 1 3
0 3
0
0 0 53616 0
4 3.3V
-12 -16 16 -8
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
972 0 0
2
43302.6 4
0
7 Ground~
168 176 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3472 0 0
2
43302.6 3
0
2 +V
167 137 100 0 1 3
0 5
0
0 0 53616 90
5 1.65V
-38 -5 -3 3
2 V2
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9998 0 0
2
43302.6 2
0
11 Signal Gen~
195 41 91 0 64 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 1070805811 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 1000 1.65 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
10 650m/2.65V
-35 -30 35 -22
2 V3
-7 -40 7 -32
0
0
39 %D %1 %2 DC 0 SIN(1.65 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
3536 0 0
2
43302.6 1
0
7 Ground~
168 83 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
4597 0 0
2
43302.6 0
0
11 Resistor:A~
219 120 86 0 2 5
0 4 7
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3835 0 0
2
43302.6 7
0
11 Resistor:A~
219 176 29 0 2 5
0 7 6
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3670 0 0
2
43302.6 6
0
8
1 3 3 0 0 4224 0 2 1 0 0 2
176 73
176 79
1 2 2 0 0 4240 0 6 5 0 0 3
83 112
83 96
72 96
1 1 4 0 0 4240 0 5 7 0 0 2
72 86
102 86
1 1 5 0 0 4240 0 4 1 0 0 2
148 98
158 98
1 4 2 0 0 16 0 3 1 0 0 2
176 112
176 105
2 5 6 0 0 8336 0 8 1 0 0 4
194 29
227 29
227 92
194 92
1 0 7 0 0 8336 0 8 0 0 8 3
158 29
146 29
146 86
2 2 7 0 0 16 0 7 1 0 0 2
138 86
158 86
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
