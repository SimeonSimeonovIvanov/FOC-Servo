CircuitMaker Text
5.6
Probes: 1
U1B_7
Transient Analysis
0 437 74 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 0 2 1
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
18
2 +V
167 293 100 0 1 3
0 5
0
0 0 53616 90
5 3.30V
-16 5 19 13
2 V7
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8396 0 0
2
5.89855e-315 0
0
11 Signal Gen~
195 36 165 0 64 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 1000 0 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 -1/1V
-18 -30 17 -22
2 V6
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(0 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3685 0 0
2
5.89855e-315 0
0
2 +V
167 293 88 0 1 3
0 6
0
0 0 53616 90
5 1.65V
-15 -16 20 -8
2 V5
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7849 0 0
2
5.89855e-315 0
0
7 Ground~
168 386 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6343 0 0
2
5.89855e-315 5.30499e-315
0
2 +V
167 386 64 0 1 3
0 7
0
0 0 53616 0
4 3.3V
-12 -16 16 -8
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7376 0 0
2
5.89855e-315 5.26354e-315
0
8 Op-Amp5~
219 386 92 0 5 11
0 3 9 7 2 8
0
0 0 848 0
10 LM6132A/NS
8 6 78 14
3 U1B
9 -14 30 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
9156 0 0
2
5.89855e-315 0
0
8 Op-Amp5~
219 176 92 0 5 11
0 12 14 10 2 13
0
0 0 848 0
10 LM6132A/NS
8 6 78 14
3 U1A
9 -14 30 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 83045552
88 0 0 256 2 1 1 0
1 U
5776 0 0
2
5.89855e-315 0
0
2 +V
167 176 64 0 1 3
0 10
0
0 0 53616 0
4 3.3V
-12 -16 16 -8
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7207 0 0
2
5.89855e-315 5.26354e-315
0
7 Ground~
168 176 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4459 0 0
2
5.89855e-315 5.30499e-315
0
2 +V
167 137 100 0 1 3
0 12
0
0 0 53616 90
5 1.65V
-38 -5 -3 3
2 V2
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3760 0 0
2
5.89855e-315 5.32571e-315
0
11 Signal Gen~
195 36 91 0 64 64
0 11 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 1070805811 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 1000 1.65 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
10 650m/2.65V
-35 -30 35 -22
2 V3
-7 -40 7 -32
0
0
39 %D %1 %2 DC 0 SIN(1.65 1 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
754 0 0
2
5.89855e-315 5.34643e-315
0
7 Ground~
168 81 186 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9767 0 0
2
5.89855e-315 5.3568e-315
0
11 Resistor:A~
219 330 160 0 2 5
0 4 3
0
0 0 880 0
2 5k
-11 20 3 28
2 R6
-12 8 2 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7978 0 0
2
5.89855e-315 0
0
11 Resistor:A~
219 330 98 0 3 5
0 5 3 1
0
0 0 880 0
2 5k
-11 20 3 28
2 R5
-12 8 2 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3142 0 0
2
5.89855e-315 0
0
11 Resistor:A~
219 386 29 0 2 5
0 9 8
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3284 0 0
2
5.89855e-315 5.30499e-315
0
11 Resistor:A~
219 330 86 0 3 5
0 6 9 1
0
0 0 880 0
2 5k
-12 -15 2 -7
2 R3
-11 -26 3 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
659 0 0
2
5.89855e-315 5.26354e-315
0
11 Resistor:A~
219 120 86 0 2 5
0 11 14
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3800 0 0
2
5.89855e-315 5.36716e-315
0
11 Resistor:A~
219 176 29 0 2 5
0 14 13
0
0 0 880 0
2 1k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6792 0 0
2
5.89855e-315 5.37752e-315
0
19
2 0 3 0 0 4096 0 14 0 0 5 2
348 98
356 98
1 1 4 0 0 4224 0 2 13 0 0 2
67 160
312 160
2 0 2 0 0 4096 0 2 0 0 13 2
67 170
81 170
1 1 5 0 0 4224 0 1 14 0 0 2
304 98
312 98
2 1 3 0 0 8320 0 13 6 0 0 4
348 160
356 160
356 98
368 98
1 1 6 0 0 4224 0 3 16 0 0 2
304 86
312 86
1 3 7 0 0 4224 0 5 6 0 0 2
386 73
386 79
1 4 2 0 0 0 0 4 6 0 0 2
386 112
386 105
2 5 8 0 0 8320 0 15 6 0 0 4
404 29
437 29
437 92
404 92
1 0 9 0 0 8320 0 15 0 0 11 3
368 29
356 29
356 86
2 2 9 0 0 0 0 16 6 0 0 2
348 86
368 86
1 3 10 0 0 4224 0 8 7 0 0 2
176 73
176 79
1 2 2 0 0 4224 0 12 11 0 0 3
81 180
81 96
67 96
1 1 11 0 0 4224 0 11 17 0 0 2
67 86
102 86
1 1 12 0 0 4224 0 10 7 0 0 2
148 98
158 98
1 4 2 0 0 0 0 9 7 0 0 2
176 112
176 105
2 5 13 0 0 8320 0 18 7 0 0 4
194 29
227 29
227 92
194 92
1 0 14 0 0 8320 0 18 0 0 19 3
158 29
146 29
146 86
2 2 14 0 0 0 0 17 7 0 0 2
138 86
158 86
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
