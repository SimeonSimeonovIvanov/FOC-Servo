CircuitMaker Text
5.6
Probes: 1
R8_2
Transient Analysis
0 473 331 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
10 10 30 100 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
2 

2 

0
0
0
39
2 +V
167 576 78 0 1 3
0 6
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3372 0 0
2
43533.5 6
0
7 Ground~
168 576 166 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3741 0 0
2
43533.5 5
0
7 Ground~
168 813 170 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5813 0 0
2
43533.5 4
0
10 Capacitor~
219 675 114 0 2 5
0 7 8
0
0 0 848 0
3 2uF
-11 -18 10 -10
2 C9
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
3213 0 0
2
43533.5 3
0
8 Coil 3T~
219 740 114 0 2 5
0 8 5
0
0 0 848 0
5 100uH
-18 -16 17 -8
2 L1
-7 -26 7 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 0 0 0 0
1 L
3694 0 0
2
43533.5 2
0
8 Op-Amp5~
219 576 114 0 5 11
0 4 7 6 2 7
0
0 0 848 0
6 OPAMP5
16 -25 58 -17
2 U3
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 0 0 0 0
1 U
4327 0 0
2
43533.5 1
0
7 Ground~
168 414 175 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8800 0 0
2
5.89823e-315 5.45523e-315
0
2 +V
167 386 157 0 1 3
0 19
0
0 0 54128 90
5 1.65V
-41 2 -6 10
2 V3
-31 -8 -17 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3406 0 0
2
5.89823e-315 5.45264e-315
0
10 Capacitor~
219 421 39 0 2 5
0 21 4
0
0 0 848 0
6 0.15nF
-22 -18 20 -10
2 C5
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6455 0 0
2
5.89823e-315 5.45005e-315
0
8 Op-Amp5~
219 414 149 0 5 11
0 19 21 22 2 4
0
0 0 848 0
7 TCA0372
5 -18 54 -10
3 U1A
19 -28 40 -20
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP16
16

0 9 10 1 13 16 9 10 1 13
16 8 7 1 4 2 0
88 0 0 256 2 1 3 0
1 U
9319 0 0
2
5.89823e-315 5.44746e-315
0
2 +V
167 414 116 0 1 3
0 22
0
0 0 54128 0
2 7V
-7 -13 7 -5
2 V2
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3172 0 0
2
5.89823e-315 5.44487e-315
0
10 Capacitor~
219 288 143 0 2 5
0 3 20
0
0 0 848 0
4 47nF
-16 -18 12 -10
2 C4
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
38 0 0
2
5.89823e-315 5.44228e-315
0
7 Ground~
168 74 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
376 0 0
2
5.89823e-315 5.43969e-315
0
11 Signal Gen~
195 35 148 0 64 64
0 9 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1176256512 0 1079194419
0 814313567 814313567 944879383 953267991 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 77105304
20
0 10000 0 3.3 0 1e-09 1e-09 5e-05 0.0001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
6 0/3.3V
-22 -30 20 -22
2 V1
-8 -40 6 -32
0
0
43 %D %1 %2 DC 0 PULSE(0 3.3 0 1n 1n 50u 100u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6666 0 0
2
5.89823e-315 5.4371e-315
0
7 Ground~
168 251 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9365 0 0
2
5.89823e-315 5.43451e-315
0
7 Ground~
168 192 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3251 0 0
2
5.89823e-315 5.43192e-315
0
7 Ground~
168 137 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5481 0 0
2
5.89823e-315 5.42933e-315
0
10 Capacitor~
219 251 169 0 2 5
0 2 3
0
0 0 848 90
4 22nF
12 0 40 8
2 C3
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7788 0 0
2
5.89823e-315 5.42414e-315
0
10 Capacitor~
219 192 168 0 2 5
0 2 24
0
0 0 848 90
4 22nF
12 0 40 8
2 C2
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3273 0 0
2
5.89823e-315 5.41896e-315
0
10 Capacitor~
219 137 167 0 2 5
0 2 23
0
0 0 848 90
4 22nF
12 0 40 8
2 C1
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3761 0 0
2
5.89823e-315 5.41378e-315
0
2 +V
167 190 409 0 1 3
0 10
0
0 0 54128 90
3 -7V
-34 2 -13 10
2 V6
-31 -8 -17 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3226 0 0
2
5.89823e-315 5.40342e-315
0
10 Capacitor~
219 110 340 0 2 5
0 9 12
0
0 0 848 0
4 47nF
-16 -18 12 -10
2 C8
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
4244 0 0
2
5.89823e-315 5.39824e-315
0
2 +V
167 412 318 0 1 3
0 16
0
0 0 54128 0
2 7V
-7 -13 7 -5
2 V7
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5225 0 0
2
5.89823e-315 5.39306e-315
0
8 Op-Amp5~
219 412 352 0 5 11
0 11 15 16 10 14
0
0 0 848 0
7 TCA0372
5 -18 54 -10
3 U2A
19 -28 40 -20
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP16
16

0 9 10 1 13 16 9 10 1 13
16 8 7 1 4 2 0
88 0 0 256 2 1 4 0
1 U
768 0 0
2
5.89823e-315 5.38788e-315
0
10 Capacitor~
219 419 241 0 2 5
0 15 14
0
0 0 848 0
5 1.5nF
-18 -18 17 -10
2 C7
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5735 0 0
2
5.89823e-315 5.37752e-315
0
2 +V
167 195 354 0 1 3
0 11
0
0 0 54128 90
2 0V
-31 2 -17 10
2 V5
-31 -8 -17 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5881 0 0
2
5.89823e-315 5.36716e-315
0
10 Capacitor~
219 242 236 0 2 5
0 17 13
0
0 0 848 0
5 1.5nF
-18 -18 17 -10
2 C6
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3275 0 0
2
5.89823e-315 5.3568e-315
0
8 Op-Amp5~
219 235 346 0 5 11
0 11 17 18 10 13
0
0 0 848 0
7 TCA0372
5 -18 54 -10
3 U1B
19 -28 40 -20
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP16
16

0 8 7 1 4 2 9 10 1 13
16 8 7 1 4 2 0
88 0 0 256 2 2 3 0
1 U
4203 0 0
2
5.89823e-315 5.34643e-315
0
2 +V
167 235 313 0 1 3
0 18
0
0 0 54128 0
2 7V
-7 -13 7 -5
2 V4
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3440 0 0
2
5.89823e-315 5.32571e-315
0
9 Resistor~
219 780 114 0 4 5
0 5 2 0 -1
0
0 0 880 0
3 100
-10 -14 11 -6
3 R10
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9102 0 0
2
43533.5 0
0
11 Resistor:A~
219 421 79 0 2 5
0 21 4
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5586 0 0
2
5.89823e-315 5.46818e-315
0
11 Resistor:A~
219 328 143 0 2 5
0 20 21
0
0 0 880 0
2 1k
-6 -14 8 -6
2 R4
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
525 0 0
2
5.89823e-315 5.46559e-315
0
11 Resistor:A~
219 113 143 0 2 5
0 9 23
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R1
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6206 0 0
2
5.89823e-315 5.463e-315
0
11 Resistor:A~
219 221 143 0 2 5
0 24 3
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R3
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3418 0 0
2
5.89823e-315 5.46041e-315
0
11 Resistor:A~
219 165 143 0 2 5
0 23 24
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R2
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9312 0 0
2
5.89823e-315 5.45782e-315
0
11 Resistor:A~
219 243 276 0 2 5
0 17 13
0
0 0 880 0
4 100k
-12 -14 16 -6
2 R7
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7419 0 0
2
5.89823e-315 5.4086e-315
0
11 Resistor:A~
219 330 346 0 2 5
0 13 15
0
0 0 880 0
4 100k
-13 -14 15 -6
2 R9
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
472 0 0
2
5.89823e-315 5.30499e-315
0
11 Resistor:A~
219 419 281 0 2 5
0 15 14
0
0 0 880 0
4 100k
-13 -14 15 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4714 0 0
2
5.89823e-315 5.26354e-315
0
11 Resistor:A~
219 149 340 0 2 5
0 12 17
0
0 0 880 0
4 100k
-12 -14 16 -6
2 R6
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9386 0 0
2
5.89823e-315 0
0
47
0 1 3 0 0 4224 0 0 12 43 0 2
251 143
279 143
1 0 4 0 0 4224 0 6 0 0 37 2
558 120
475 120
2 1 2 0 0 8320 0 30 3 0 0 3
798 114
813 114
813 164
1 2 5 0 0 4224 0 30 5 0 0 2
762 114
760 114
1 3 6 0 0 4224 0 1 6 0 0 2
576 87
576 101
1 4 2 0 0 0 0 2 6 0 0 2
576 160
576 127
1 0 7 0 0 4096 0 4 0 0 8 2
666 114
642 114
2 5 7 0 0 12416 0 6 6 0 0 6
558 108
531 108
531 39
642 39
642 114
594 114
2 1 8 0 0 4224 0 4 5 0 0 2
684 114
720 114
1 0 9 0 0 8320 0 22 0 0 39 3
101 340
88 340
88 143
4 0 10 0 0 4096 0 28 0 0 12 2
235 359
235 407
4 1 10 0 0 8320 0 24 21 0 0 3
412 365
412 407
201 407
0 1 11 0 0 8320 0 0 24 22 0 5
211 352
211 382
362 382
362 358
394 358
2 1 12 0 0 4224 0 22 39 0 0 2
119 340
131 340
1 0 13 0 0 4096 0 37 0 0 28 2
312 346
296 346
2 0 14 0 0 4096 0 25 0 0 21 3
428 241
473 241
473 281
1 0 15 0 0 4096 0 25 0 0 18 3
410 241
365 241
365 281
1 0 15 0 0 8320 0 38 0 0 19 3
401 281
365 281
365 346
2 2 15 0 0 0 0 37 24 0 0 2
348 346
394 346
1 3 16 0 0 4224 0 23 24 0 0 2
412 327
412 339
5 2 14 0 0 8320 0 24 38 0 0 4
430 352
473 352
473 281
437 281
1 1 11 0 0 0 0 26 28 0 0 2
206 352
217 352
2 0 13 0 0 4096 0 27 0 0 28 3
251 236
296 236
296 276
1 0 17 0 0 4096 0 27 0 0 25 3
233 236
188 236
188 276
1 0 17 0 0 8320 0 36 0 0 26 3
225 276
188 276
188 340
2 2 17 0 0 0 0 39 28 0 0 2
167 340
217 340
1 3 18 0 0 4224 0 29 28 0 0 2
235 322
235 333
5 2 13 0 0 8320 0 28 36 0 0 4
253 346
296 346
296 276
261 276
1 4 2 0 0 0 0 7 10 0 0 2
414 169
414 162
1 1 19 0 0 4224 0 8 10 0 0 2
397 155
396 155
2 1 20 0 0 4224 0 12 32 0 0 2
297 143
310 143
2 0 4 0 0 0 0 9 0 0 37 3
430 39
475 39
475 79
1 0 21 0 0 4096 0 9 0 0 34 3
412 39
367 39
367 79
1 0 21 0 0 8320 0 31 0 0 35 3
403 79
367 79
367 143
2 2 21 0 0 0 0 32 10 0 0 2
346 143
396 143
1 3 22 0 0 4224 0 11 10 0 0 2
414 125
414 136
5 2 4 0 0 128 0 10 31 0 0 4
432 149
475 149
475 79
439 79
1 2 2 0 0 128 0 13 14 0 0 3
74 184
74 153
66 153
1 1 9 0 0 0 0 14 33 0 0 2
66 143
95 143
1 1 2 0 0 0 0 15 18 0 0 2
251 184
251 178
1 1 2 0 0 0 0 16 19 0 0 2
192 184
192 177
1 1 2 0 0 0 0 17 20 0 0 2
137 184
137 176
2 2 3 0 0 128 0 34 18 0 0 3
239 143
251 143
251 160
2 0 23 0 0 4096 0 20 0 0 47 2
137 158
137 143
2 0 24 0 0 4096 0 19 0 0 46 2
192 159
192 143
2 1 24 0 0 4224 0 35 34 0 0 2
183 143
203 143
2 1 23 0 0 4224 0 33 35 0 0 2
131 143
147 143
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.003 2e-07 2e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
