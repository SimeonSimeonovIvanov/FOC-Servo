CircuitMaker Text
5.6
Probes: 1
V1_1
Transient Analysis
0 90 141 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
2 

2 

0
0
0
65
10 Capacitor~
219 966 541 0 2 5
0 3 3
0
0 0 848 180
3 1uF
-11 -18 10 -10
3 C15
-11 -28 10 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
388 0 0
2
43562.7 0
0
7 Ground~
168 445 457 0 1 3
0 2
0
0 0 53360 270
0
5 GND14
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4595 0 0
2
43562.7 0
0
7 Ground~
168 446 501 0 1 3
0 2
0
0 0 53360 270
0
5 GND13
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3173 0 0
2
43562.7 0
0
7 Ground~
168 575 607 0 1 3
0 2
0
0 0 53360 0
0
5 GND12
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9261 0 0
2
43562.7 0
0
10 Capacitor~
219 501 516 0 2 5
0 5 2
0
0 0 848 90
3 1nF
18 0 39 8
3 C14
18 -10 39 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3494 0 0
2
43562.7 0
0
10 Capacitor~
219 501 485 0 2 5
0 2 6
0
0 0 848 90
3 1nF
18 0 39 8
3 C13
18 -10 39 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9101 0 0
2
43562.7 0
0
2 +V
167 614 512 0 1 3
0 10
0
0 0 54256 0
4 +15V
-15 -22 13 -14
3 V10
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
358 0 0
2
43562.7 2
0
7 Ground~
168 614 607 0 1 3
0 2
0
0 0 53360 0
0
5 GND11
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3726 0 0
2
43562.7 1
0
8 Op-Amp5~
219 614 548 0 5 11
0 9 7 10 2 8
0
0 0 848 0
6 OPAMP5
16 -25 58 -17
2 U5
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
999 0 0
2
43562.7 0
0
7 Ground~
168 924 628 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8787 0 0
2
43562.7 0
0
10 Capacitor~
219 924 605 0 2 5
0 2 11
0
0 0 848 90
4 47nF
14 0 42 8
3 C12
18 -10 39 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
3348 0 0
2
43562.7 0
0
7 Ground~
168 799 594 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3395 0 0
2
43562.7 0
0
10 Capacitor~
219 799 567 0 2 5
0 2 12
0
0 0 848 90
5 1.2nF
11 0 46 8
3 C11
18 -10 39 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7740 0 0
2
43562.7 0
0
10 Capacitor~
219 742 499 0 2 5
0 13 3
0
0 0 848 90
5 4.7nF
11 0 46 8
3 C10
18 -10 39 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6480 0 0
2
43562.7 0
0
8 Op-Amp5~
219 858 542 0 5 11
0 12 3 14 2 3
0
0 0 848 0
6 OPAMP5
16 -25 58 -17
2 U4
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
342 0 0
2
43562.7 2
0
7 Ground~
168 858 594 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9953 0 0
2
43562.7 1
0
2 +V
167 858 506 0 1 3
0 14
0
0 0 54256 0
4 +15V
-15 -22 13 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
361 0 0
2
43562.7 0
0
2 +V
167 576 78 0 1 3
0 18
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V9
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3343 0 0
2
5.89884e-315 5.36716e-315
0
7 Ground~
168 576 166 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7923 0 0
2
5.89884e-315 5.3568e-315
0
7 Ground~
168 813 170 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6174 0 0
2
5.89884e-315 5.34643e-315
0
10 Capacitor~
219 675 114 0 2 5
0 19 20
0
0 0 848 0
3 2uF
-11 -18 10 -10
2 C9
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6692 0 0
2
5.89884e-315 5.32571e-315
0
8 Coil 3T~
219 740 114 0 2 5
0 20 17
0
0 0 848 0
5 100uH
-18 -16 17 -8
2 L1
-7 -26 7 -18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
76 0 0 0 1 0 0 0
1 L
8790 0 0
2
5.89884e-315 5.30499e-315
0
8 Op-Amp5~
219 576 114 0 5 11
0 16 19 18 2 19
0
0 0 848 0
6 OPAMP5
16 -25 58 -17
2 U3
30 -35 44 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
4595 0 0
2
5.89884e-315 5.26354e-315
0
7 Ground~
168 414 175 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
667 0 0
2
43562.7 0
0
2 +V
167 386 157 0 1 3
0 30
0
0 0 54128 90
5 1.65V
-41 2 -6 10
2 V3
-31 -8 -17 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8743 0 0
2
43562.7 1
0
10 Capacitor~
219 421 39 0 2 5
0 32 16
0
0 0 848 0
6 0.15nF
-22 -18 20 -10
2 C5
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8298 0 0
2
43562.7 2
0
8 Op-Amp5~
219 414 149 0 5 11
0 30 32 33 2 16
0
0 0 848 0
7 TCA0372
5 -18 54 -10
3 U1A
19 -28 40 -20
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP16
16

0 9 10 1 13 16 9 10 1 13
16 8 7 1 4 2 0
88 0 0 256 2 1 3 0
1 U
313 0 0
2
43562.7 3
0
2 +V
167 414 116 0 1 3
0 33
0
0 0 54128 0
2 7V
-7 -13 7 -5
2 V2
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7548 0 0
2
43562.7 4
0
10 Capacitor~
219 288 143 0 2 5
0 15 31
0
0 0 848 0
4 47nF
-16 -18 12 -10
2 C4
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8973 0 0
2
43562.7 5
0
7 Ground~
168 74 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9712 0 0
2
43562.7 6
0
11 Signal Gen~
195 35 148 0 64 64
0 4 2 1 86 -10 10 0 0 0
0 0 0 0 0 0 0 1176256512 0 1079194419
0 814313567 814313567 944879383 953267991 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 77105304
20
0 10000 0 3.3 0 1e-09 1e-09 5e-05 0.0001 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
6 0/3.3V
-22 -30 20 -22
2 V1
-8 -40 6 -32
0
0
43 %D %1 %2 DC 0 PULSE(0 3.3 0 1n 1n 50u 100u)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4518 0 0
2
43562.7 7
0
7 Ground~
168 251 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5596 0 0
2
43562.7 8
0
7 Ground~
168 192 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
692 0 0
2
43562.7 9
0
7 Ground~
168 137 190 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6258 0 0
2
43562.7 10
0
10 Capacitor~
219 251 169 0 2 5
0 2 15
0
0 0 848 90
4 22nF
12 0 40 8
2 C3
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5578 0 0
2
43562.7 11
0
10 Capacitor~
219 192 168 0 2 5
0 2 35
0
0 0 848 90
4 22nF
12 0 40 8
2 C2
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
8709 0 0
2
43562.7 12
0
10 Capacitor~
219 137 167 0 2 5
0 2 34
0
0 0 848 90
4 22nF
12 0 40 8
2 C1
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
9131 0 0
2
43562.7 13
0
2 +V
167 190 409 0 1 3
0 21
0
0 0 54128 90
3 -7V
-34 2 -13 10
2 V6
-31 -8 -17 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3645 0 0
2
43562.7 14
0
10 Capacitor~
219 110 340 0 2 5
0 4 23
0
0 0 848 0
4 47nF
-16 -18 12 -10
2 C8
-9 -28 5 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7613 0 0
2
43562.7 15
0
2 +V
167 412 318 0 1 3
0 27
0
0 0 54128 0
2 7V
-7 -13 7 -5
2 V7
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9467 0 0
2
43562.7 16
0
8 Op-Amp5~
219 412 352 0 5 11
0 22 26 27 21 25
0
0 0 848 0
7 TCA0372
5 -18 54 -10
3 U2A
19 -28 40 -20
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP16
16

0 9 10 1 13 16 9 10 1 13
16 8 7 1 4 2 0
88 0 0 256 2 1 4 0
1 U
3932 0 0
2
43562.7 17
0
10 Capacitor~
219 419 241 0 2 5
0 26 25
0
0 0 848 0
5 1.5nF
-18 -18 17 -10
2 C7
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5288 0 0
2
43562.7 18
0
2 +V
167 195 354 0 1 3
0 22
0
0 0 54128 90
2 0V
-31 2 -17 10
2 V5
-31 -8 -17 0
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4934 0 0
2
43562.7 19
0
10 Capacitor~
219 242 236 0 2 5
0 28 24
0
0 0 848 0
5 1.5nF
-18 -18 17 -10
2 C6
-8 -28 6 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
5987 0 0
2
43562.7 20
0
8 Op-Amp5~
219 235 346 0 5 11
0 22 28 29 21 24
0
0 0 848 0
7 TCA0372
5 -18 54 -10
3 U1B
19 -28 40 -20
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 DIP16
16

0 8 7 1 4 2 9 10 1 13
16 8 7 1 4 2 0
88 0 0 256 2 2 3 0
1 U
7737 0 0
2
43562.7 21
0
2 +V
167 235 313 0 1 3
0 29
0
0 0 54128 0
2 7V
-7 -13 7 -5
2 V4
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4200 0 0
2
43562.7 22
0
11 Resistor:A~
219 475 458 0 3 5
0 2 6 -1
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R19
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5780 0 0
2
43562.7 0
0
11 Resistor:A~
219 473 554 0 2 5
0 4 5
0
0 0 880 0
3 10k
-10 -14 11 -6
3 R18
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6490 0 0
2
43562.7 0
0
11 Resistor:A~
219 541 458 0 2 5
0 6 7
0
0 0 880 0
4 5.1k
-13 -14 15 -6
3 R17
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8663 0 0
2
43562.7 0
0
11 Resistor:A~
219 541 554 0 2 5
0 5 9
0
0 0 880 0
4 5.1k
-13 -14 15 -6
3 R16
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
318 0 0
2
43562.7 0
0
11 Resistor:A~
219 575 579 0 3 5
0 2 9 -1
0
0 0 880 90
3 68k
12 0 33 8
3 R15
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
348 0 0
2
43562.7 0
0
11 Resistor:A~
219 613 458 0 2 5
0 7 8
0
0 0 880 0
3 68k
-10 -14 11 -6
3 R14
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8551 0 0
2
43562.7 0
0
11 Resistor:A~
219 924 570 0 2 5
0 11 3
0
0 0 880 90
2 47
15 0 29 8
3 R13
11 -10 32 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7295 0 0
2
43562.7 0
0
11 Resistor:A~
219 714 548 0 2 5
0 8 13
0
0 0 880 0
4 3.3k
-13 -14 15 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9900 0 0
2
43562.7 0
0
11 Resistor:A~
219 769 548 0 2 5
0 13 12
0
0 0 880 0
4 3.3k
-13 -14 15 -6
3 R11
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8725 0 0
2
43562.7 0
0
9 Resistor~
219 780 114 0 4 5
0 17 2 0 -1
0
0 0 880 0
3 100
-10 -14 11 -6
3 R10
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
366 0 0
2
5.89884e-315 0
0
11 Resistor:A~
219 421 79 0 2 5
0 32 16
0
0 0 880 0
3 10k
-10 -14 11 -6
2 R5
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5762 0 0
2
43562.7 23
0
11 Resistor:A~
219 328 143 0 2 5
0 31 32
0
0 0 880 0
2 1k
-6 -14 8 -6
2 R4
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4943 0 0
2
43562.7 24
0
11 Resistor:A~
219 113 143 0 2 5
0 4 34
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R1
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3435 0 0
2
43562.7 25
0
11 Resistor:A~
219 221 143 0 2 5
0 35 15
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R3
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8705 0 0
2
43562.7 26
0
11 Resistor:A~
219 165 143 0 2 5
0 34 35
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R2
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4331 0 0
2
43562.7 27
0
11 Resistor:A~
219 243 276 0 2 5
0 28 24
0
0 0 880 0
4 100k
-12 -14 16 -6
2 R7
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
787 0 0
2
43562.7 28
0
11 Resistor:A~
219 330 346 0 2 5
0 24 26
0
0 0 880 0
4 100k
-13 -14 15 -6
2 R9
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3655 0 0
2
43562.7 29
0
11 Resistor:A~
219 419 281 0 2 5
0 26 25
0
0 0 880 0
4 100k
-13 -14 15 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6682 0 0
2
43562.7 30
0
11 Resistor:A~
219 149 340 0 2 5
0 23 28
0
0 0 880 0
4 100k
-12 -14 16 -6
2 R6
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
582 0 0
2
43562.7 31
0
78
1 0 3 0 0 12288 0 1 0 0 2 5
975 541
991 541
991 560
944 560
944 541
0 2 3 0 0 0 0 0 1 22 0 3
924 542
924 541
957 541
1 0 4 0 0 4224 0 48 0 0 41 3
455 554
88 554
88 340
1 1 2 0 0 4096 0 2 47 0 0 2
452 458
457 458
2 0 5 0 0 4096 0 48 0 0 9 2
491 554
501 554
2 0 6 0 0 4096 0 47 0 0 10 2
493 458
501 458
1 0 2 0 0 4096 0 3 0 0 11 2
453 502
501 502
1 1 2 0 0 0 0 4 51 0 0 2
575 601
575 597
1 1 5 0 0 8320 0 50 5 0 0 3
523 554
501 554
501 525
1 2 6 0 0 4224 0 49 6 0 0 3
523 458
501 458
501 476
2 1 2 0 0 0 0 5 6 0 0 2
501 507
501 494
2 0 7 0 0 4096 0 49 0 0 14 2
559 458
575 458
2 0 8 0 0 8320 0 52 0 0 17 3
631 458
673 458
673 548
2 1 7 0 0 8320 0 9 52 0 0 4
596 542
575 542
575 458
595 458
2 0 9 0 0 4096 0 51 0 0 16 2
575 561
575 554
2 1 9 0 0 4224 0 50 9 0 0 2
559 554
596 554
5 1 8 0 0 0 0 9 54 0 0 2
632 548
696 548
1 3 10 0 0 4224 0 7 9 0 0 2
614 521
614 535
1 4 2 0 0 0 0 8 9 0 0 2
614 601
614 561
1 1 2 0 0 0 0 10 11 0 0 2
924 622
924 614
2 1 11 0 0 4224 0 11 53 0 0 2
924 596
924 588
2 0 3 0 0 0 0 53 0 0 29 2
924 552
924 542
2 0 12 0 0 4096 0 13 0 0 28 2
799 558
799 548
1 1 2 0 0 0 0 12 13 0 0 2
799 588
799 576
2 0 3 0 0 8192 0 14 0 0 29 3
742 490
742 458
824 458
1 0 13 0 0 4224 0 14 0 0 27 2
742 508
742 548
2 1 13 0 0 0 0 54 55 0 0 2
732 548
751 548
2 1 12 0 0 4224 0 55 15 0 0 2
787 548
840 548
2 5 3 0 0 12416 0 15 15 0 0 6
840 536
824 536
824 458
924 458
924 542
876 542
1 3 14 0 0 4224 0 17 15 0 0 2
858 515
858 529
1 4 2 0 0 0 0 16 15 0 0 2
858 588
858 555
0 1 15 0 0 4224 0 0 29 74 0 2
251 143
279 143
1 0 16 0 0 4224 0 23 0 0 68 2
558 120
475 120
2 1 2 0 0 8320 0 56 20 0 0 3
798 114
813 114
813 164
1 2 17 0 0 4224 0 56 22 0 0 2
762 114
760 114
1 3 18 0 0 4224 0 18 23 0 0 2
576 87
576 101
1 4 2 0 0 0 0 19 23 0 0 2
576 160
576 127
1 0 19 0 0 4096 0 21 0 0 39 2
666 114
642 114
2 5 19 0 0 12416 0 23 23 0 0 6
558 108
531 108
531 39
642 39
642 114
594 114
2 1 20 0 0 4224 0 21 22 0 0 2
684 114
720 114
1 0 4 0 0 128 0 39 0 0 70 3
101 340
88 340
88 143
4 0 21 0 0 4096 0 45 0 0 43 2
235 359
235 407
4 1 21 0 0 8320 0 41 38 0 0 3
412 365
412 407
201 407
0 1 22 0 0 8320 0 0 41 53 0 5
211 352
211 382
362 382
362 358
394 358
2 1 23 0 0 4224 0 39 65 0 0 2
119 340
131 340
1 0 24 0 0 4096 0 63 0 0 59 2
312 346
296 346
2 0 25 0 0 4096 0 42 0 0 52 3
428 241
473 241
473 281
1 0 26 0 0 4096 0 42 0 0 49 3
410 241
365 241
365 281
1 0 26 0 0 8320 0 64 0 0 50 3
401 281
365 281
365 346
2 2 26 0 0 0 0 63 41 0 0 2
348 346
394 346
1 3 27 0 0 4224 0 40 41 0 0 2
412 327
412 339
5 2 25 0 0 8320 0 41 64 0 0 4
430 352
473 352
473 281
437 281
1 1 22 0 0 0 0 43 45 0 0 2
206 352
217 352
2 0 24 0 0 4096 0 44 0 0 59 3
251 236
296 236
296 276
1 0 28 0 0 4096 0 44 0 0 56 3
233 236
188 236
188 276
1 0 28 0 0 8320 0 62 0 0 57 3
225 276
188 276
188 340
2 2 28 0 0 0 0 65 45 0 0 2
167 340
217 340
1 3 29 0 0 4224 0 46 45 0 0 2
235 322
235 333
5 2 24 0 0 8320 0 45 62 0 0 4
253 346
296 346
296 276
261 276
1 4 2 0 0 0 0 24 27 0 0 2
414 169
414 162
1 1 30 0 0 4224 0 25 27 0 0 2
397 155
396 155
2 1 31 0 0 4224 0 29 58 0 0 2
297 143
310 143
2 0 16 0 0 0 0 26 0 0 68 3
430 39
475 39
475 79
1 0 32 0 0 4096 0 26 0 0 65 3
412 39
367 39
367 79
1 0 32 0 0 8320 0 57 0 0 66 3
403 79
367 79
367 143
2 2 32 0 0 0 0 58 27 0 0 2
346 143
396 143
1 3 33 0 0 4224 0 28 27 0 0 2
414 125
414 136
5 2 16 0 0 0 0 27 57 0 0 4
432 149
475 149
475 79
439 79
1 2 2 0 0 0 0 30 31 0 0 3
74 184
74 153
66 153
1 1 4 0 0 0 0 31 59 0 0 2
66 143
95 143
1 1 2 0 0 0 0 32 35 0 0 2
251 184
251 178
1 1 2 0 0 0 0 33 36 0 0 2
192 184
192 177
1 1 2 0 0 0 0 34 37 0 0 2
137 184
137 176
2 2 15 0 0 0 0 60 35 0 0 3
239 143
251 143
251 160
2 0 34 0 0 4096 0 37 0 0 78 2
137 158
137 143
2 0 35 0 0 4096 0 36 0 0 77 2
192 159
192 143
2 1 35 0 0 4224 0 61 60 0 0 2
183 143
203 143
2 1 34 0 0 4224 0 59 61 0 0 2
131 143
147 143
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-07 2e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
