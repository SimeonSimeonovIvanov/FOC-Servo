CircuitMaker Text
5.6
Probes: 1
U1B_7
Transient Analysis
0 665 109 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 240 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
20
8 Op-Amp5~
219 638 111 0 5 11
0 8 9 10 2 11
0
0 0 848 0
5 LM358
11 6 46 14
3 U1B
12 -13 33 -5
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
6901 0 0
2
43544 0
0
2 +V
167 591 185 0 1 3
0 7
0
0 0 54128 180
1 0
-2 12 5 20
5 Vref2
-15 1 20 9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
842 0 0
2
43544 1
0
11 Signal Gen~
195 399 112 0 64 64
0 5 6 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846080 1075838976 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 1000 2.5 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 2/3V
-15 -30 13 -22
2 V4
-8 -40 6 -32
0
0
34 %D %1 %2 DC 0 SIN(2.5 500m 1k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3277 0 0
2
43544 2
0
7 Ground~
168 638 137 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4212 0 0
2
43544 3
0
2 +V
167 638 78 0 1 3
0 10
0
0 0 54128 0
2 10
-6 -13 8 -5
2 V3
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4720 0 0
2
43544 4
0
2 +V
167 287 69 0 1 3
0 15
0
0 0 54128 0
2 10
-6 -13 8 -5
2 V2
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5551 0 0
2
43544 5
0
7 Ground~
168 287 128 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6986 0 0
2
43544 6
0
11 Signal Gen~
195 48 103 0 64 64
0 3 4 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846080 0 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 1000 0 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -500m/500mV
-39 -30 38 -22
2 V1
-8 -40 6 -32
0
0
32 %D %1 %2 DC 0 SIN(0 500m 1k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8745 0 0
2
43544 7
0
2 +V
167 240 176 0 1 3
0 12
0
0 0 54128 180
4 1.65
-12 12 16 20
5 Vref1
-15 1 20 9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9592 0 0
2
43544 8
0
8 Op-Amp5~
219 287 102 0 5 11
0 13 14 15 2 16
0
0 0 848 0
5 LM358
11 6 46 14
3 U1A
12 -13 33 -5
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
8748 0 0
2
43544 9
0
11 Resistor:A~
219 500 112 0 2 5
0 5 6
0
0 0 880 90
3 120
7 0 28 8
3 R10
8 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
43544 10
0
11 Resistor:A~
219 552 117 0 2 5
0 5 8
0
0 0 880 0
2 3k
-6 16 8 24
2 R9
-11 6 3 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
631 0 0
2
43544 11
0
11 Resistor:A~
219 591 147 0 3 5
0 7 8 1
0
0 0 880 90
2 3k
10 0 24 8
2 R8
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9466 0 0
2
43544 12
0
11 Resistor:A~
219 552 105 0 2 5
0 6 9
0
0 0 880 0
2 3k
-6 -14 8 -6
2 R5
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3266 0 0
2
43544 13
0
11 Resistor:A~
219 635 41 0 2 5
0 9 11
0
0 0 880 0
2 3k
-6 -14 8 -6
2 R4
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7693 0 0
2
43544 14
0
11 Resistor:A~
219 284 32 0 2 5
0 14 16
0
0 0 880 0
2 3k
-6 -14 8 -6
2 R7
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3723 0 0
2
43544 15
0
11 Resistor:A~
219 201 96 0 2 5
0 4 14
0
0 0 880 0
2 3k
-6 -14 8 -6
2 R6
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3440 0 0
2
43544 16
0
11 Resistor:A~
219 240 138 0 3 5
0 12 13 1
0
0 0 880 90
2 3k
10 0 24 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6263 0 0
2
43544 17
0
11 Resistor:A~
219 201 108 0 2 5
0 3 13
0
0 0 880 0
2 3k
-6 16 8 24
2 R2
-11 6 3 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4900 0 0
2
43544 18
0
11 Resistor:A~
219 149 103 0 2 5
0 3 4
0
0 0 880 90
3 120
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8783 0 0
2
43544 19
0
24
1 0 3 0 0 12416 0 8 0 0 17 4
79 98
97 98
97 126
150 126
2 0 4 0 0 12416 0 8 0 0 16 4
79 108
111 108
111 78
149 78
1 0 5 0 0 12416 0 3 0 0 7 4
430 107
448 107
448 135
500 135
2 0 6 0 0 12416 0 3 0 0 6 4
430 117
463 117
463 87
500 87
1 1 7 0 0 4224 0 2 13 0 0 2
591 170
591 165
2 1 6 0 0 0 0 11 14 0 0 5
500 94
500 87
528 87
528 105
534 105
1 1 5 0 0 0 0 12 11 0 0 5
534 117
528 117
528 135
500 135
500 130
2 0 8 0 0 4096 0 13 0 0 9 2
591 129
591 117
2 1 8 0 0 4224 0 12 1 0 0 2
570 117
620 117
1 4 2 0 0 4224 0 4 1 0 0 2
638 131
638 124
1 0 9 0 0 8320 0 15 0 0 12 3
617 41
591 41
591 105
2 2 9 0 0 0 0 14 1 0 0 2
570 105
620 105
1 3 10 0 0 4224 0 5 1 0 0 2
638 87
638 98
5 2 11 0 0 8320 0 1 15 0 0 4
656 111
683 111
683 41
653 41
1 1 12 0 0 4224 0 9 18 0 0 2
240 161
240 156
2 1 4 0 0 0 0 20 17 0 0 5
149 85
149 78
177 78
177 96
183 96
1 1 3 0 0 0 0 19 20 0 0 5
183 108
177 108
177 126
149 126
149 121
2 0 13 0 0 4096 0 18 0 0 19 2
240 120
240 108
2 1 13 0 0 4224 0 19 10 0 0 2
219 108
269 108
1 4 2 0 0 0 0 7 10 0 0 2
287 122
287 115
1 0 14 0 0 8320 0 16 0 0 22 3
266 32
240 32
240 96
2 2 14 0 0 0 0 17 10 0 0 2
219 96
269 96
1 3 15 0 0 4224 0 6 10 0 0 2
287 78
287 89
5 2 16 0 0 8320 0 10 16 0 0 4
305 102
332 102
332 32
302 32
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
