CircuitMaker Text
5.6
Probes: 1
R12_2
Transient Analysis
0 642 97 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 170 10
445 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.410638 0.500000
613 175 1743 561
9961490 0
0
6 Title:
5 Name:
0
0
0
32
11 Signal Gen~
195 426 98 0 64 64
0 4 3 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1120403456 0 1092616192
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 264
20
1 100 0 10 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -10/10V
-25 -30 24 -22
2 V5
-8 -40 6 -32
0
0
38 %D %1 %2 DC 0 SIN(0 10 100 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4316 0 0
2
43325.9 0
0
8 Op-Amp5~
219 621 98 0 5 11
0 12 13 16 2 15
0
0 0 848 0
6 OP284E
11 6 53 14
3 U2B
9 -14 30 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 2 0
1 U
3315 0 0
2
43325.8 0
0
2 +V
167 473 301 0 1 3
0 7
0
0 0 53616 90
2 0V
-21 -6 -7 2
2 V8
-43 -15 -29 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7100 0 0
2
43325.8 1
0
11 Signal Gen~
195 425 235 0 64 64
0 5 3 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1120403456 1084227584 1084227584
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 40691264
20
1 100 5 5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
5 0/10V
-19 -30 16 -22
2 V6
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(5 5 100 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8968 0 0
2
43325.8 0
0
8 Op-Amp5~
219 595 246 0 5 11
0 8 9 11 2 10
0
0 0 848 0
6 OP284E
11 7 53 15
3 U2A
9 -17 30 -9
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 110
88 0 0 256 2 1 2 0
1 U
3557 0 0
2
43325.8 0
0
2 +V
167 595 211 0 1 3
0 11
0
0 0 53616 0
4 3.3V
-13 -16 15 -8
2 V7
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6695 0 0
2
43325.8 4
0
7 Ground~
168 595 280 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5921 0 0
2
43325.8 3
0
2 +V
167 492 147 0 1 3
0 14
0
0 0 53616 90
5 1.65V
-40 -6 -5 2
3 V11
-46 -15 -25 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3726 0 0
2
5.89855e-315 5.32571e-315
0
7 Ground~
168 621 132 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6207 0 0
2
5.89855e-315 5.26354e-315
0
2 +V
167 621 63 0 1 3
0 16
0
0 0 53616 0
4 3.3V
-13 -16 15 -8
3 V13
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7606 0 0
2
5.89855e-315 0
0
7 Ground~
168 69 156 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
915 0 0
2
5.89855e-315 0
0
11 Signal Gen~
195 30 103 0 64 64
0 18 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1092616192
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 70
20
1 1000 0 10 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -10/10V
-25 -30 24 -22
2 V4
-8 -40 6 -32
0
0
37 %D %1 %2 DC 0 SIN(0 10 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5257 0 0
2
5.89855e-315 5.26354e-315
0
7 Ground~
168 129 156 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7821 0 0
2
5.89855e-315 5.30499e-315
0
2 +V
167 206 141 0 1 3
0 19
0
0 0 54128 90
5 3.30V
-39 -5 -4 3
2 V3
-29 -15 -15 -7
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3906 0 0
2
5.89855e-315 5.32571e-315
0
2 +V
167 210 88 0 1 3
0 21
0
0 0 54128 90
5 1.65V
-38 -6 -3 2
2 V2
-28 -16 -14 -8
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9214 0 0
2
5.89855e-315 5.34643e-315
0
7 Ground~
168 303 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6348 0 0
2
5.89855e-315 5.3568e-315
0
2 +V
167 303 64 0 1 3
0 22
0
0 0 54128 0
4 3.3V
-12 -16 16 -8
2 V1
-5 -26 9 -18
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6354 0 0
2
5.89855e-315 5.36716e-315
0
8 Op-Amp5~
219 303 92 0 5 11
0 20 24 22 2 23
0
0 0 848 0
10 LM6132A/NS
8 6 78 14
3 U1B
9 -14 30 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
4426 0 0
2
5.89855e-315 5.37752e-315
0
11 Resistor:A~
219 528 299 0 3 5
0 7 8 1
0
0 0 880 0
3 10k
-9 21 12 29
2 R7
-6 8 8 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9745 0 0
2
43325.8 0
0
11 Resistor:A~
219 527 252 0 2 5
0 5 8
0
0 0 880 0
3 33k
-10 16 11 24
3 R16
-10 6 11 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4804 0 0
2
43325.8 9
0
11 Resistor:A~
219 527 240 0 2 5
0 3 9
0
0 0 880 0
3 33k
-10 -14 11 -6
3 R15
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8371 0 0
2
43325.8 8
0
11 Resistor:A~
219 558 216 0 2 5
0 9 10
0
0 0 880 90
3 10k
4 0 25 8
2 R9
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
697 0 0
2
43325.8 7
0
11 Resistor:A~
219 552 145 0 3 5
0 14 12 1
0
0 0 880 0
4 5.1k
-13 21 15 29
3 R10
-9 8 12 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3889 0 0
2
5.89855e-315 5.39306e-315
0
11 Resistor:A~
219 584 68 0 2 5
0 13 15
0
0 0 880 90
4 5.1k
6 0 34 8
3 R12
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6643 0 0
2
5.89855e-315 5.37752e-315
0
11 Resistor:A~
219 553 92 0 2 5
0 4 13
0
0 0 880 0
3 33k
-10 -14 11 -6
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8554 0 0
2
5.89855e-315 5.36716e-315
0
11 Resistor:A~
219 553 104 0 2 5
0 3 12
0
0 0 880 0
3 33k
-10 16 11 24
3 R14
-10 6 11 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9989 0 0
2
5.89855e-315 5.3568e-315
0
11 Resistor:A~
219 103 98 0 2 5
0 18 17
0
0 0 880 0
4 6.2k
-12 8 16 16
2 R6
-11 -14 3 -6
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3137 0 0
2
5.89855e-315 5.38788e-315
0
11 Resistor:A~
219 129 124 0 3 5
0 2 17 -1
0
0 0 880 90
4 1.1k
8 0 36 8
2 R5
15 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7969 0 0
2
5.89855e-315 5.39306e-315
0
11 Resistor:A~
219 246 139 0 3 5
0 19 20 1
0
0 0 880 0
3 51k
-14 20 7 28
2 R4
-11 10 3 18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5719 0 0
2
5.89855e-315 5.39824e-315
0
11 Resistor:A~
219 247 98 0 2 5
0 17 20
0
0 0 880 0
3 51k
-14 20 7 28
2 R3
-11 10 3 18
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5243 0 0
2
5.89855e-315 5.40342e-315
0
11 Resistor:A~
219 303 29 0 2 5
0 24 23
0
0 0 880 0
3 51k
-10 -14 11 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8250 0 0
2
5.89855e-315 5.4086e-315
0
11 Resistor:A~
219 247 86 0 3 5
0 21 24 1
0
0 0 880 0
3 51k
-15 -15 6 -7
2 R1
-12 -25 2 -17
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8570 0 0
2
5.89855e-315 5.41378e-315
0
36
0 0 3 0 0 12432 0 0 0 2 5 6
468 103
468 131
371 131
371 277
467 277
467 240
2 1 3 0 0 128 0 1 26 0 0 4
457 103
520 103
520 104
535 104
1 1 4 0 0 4224 0 1 25 0 0 4
457 93
520 93
520 92
535 92
1 1 5 0 0 4224 0 4 20 0 0 4
456 230
489 230
489 252
509 252
1 2 3 0 0 128 0 21 4 0 0 2
509 240
456 240
0 0 6 0 0 128 0 0 0 0 0 2
558 353
558 353
1 1 7 0 0 4224 0 3 19 0 0 2
484 299
510 299
0 2 8 0 0 4224 0 0 19 10 0 3
558 252
558 299
546 299
1 0 9 0 0 4096 0 22 0 0 12 2
558 234
558 240
2 1 8 0 0 128 0 20 5 0 0 2
545 252
577 252
2 5 10 0 0 8320 0 22 5 0 0 5
558 198
558 186
672 186
672 246
613 246
2 2 9 0 0 4224 0 21 5 0 0 2
545 240
577 240
1 4 2 0 0 4096 0 7 5 0 0 2
595 274
595 259
3 1 11 0 0 4224 0 5 6 0 0 2
595 233
595 220
2 0 12 0 0 8320 0 23 0 0 17 3
570 145
584 145
584 104
1 0 13 0 0 4096 0 24 0 0 20 2
584 86
584 92
2 1 12 0 0 0 0 26 2 0 0 2
571 104
603 104
1 1 14 0 0 4224 0 8 23 0 0 2
503 145
534 145
2 5 15 0 0 8320 0 24 2 0 0 5
584 50
584 38
672 38
672 98
639 98
2 2 13 0 0 4224 0 25 2 0 0 2
571 92
603 92
1 4 2 0 0 0 0 9 2 0 0 2
621 126
621 111
3 1 16 0 0 4224 0 2 10 0 0 2
621 85
621 72
1 0 17 0 0 4224 0 30 0 0 27 2
229 98
129 98
1 1 18 0 0 4224 0 12 27 0 0 2
61 98
85 98
1 2 2 0 0 4224 0 11 12 0 0 3
69 150
69 108
61 108
1 1 2 0 0 0 0 13 28 0 0 2
129 150
129 142
2 2 17 0 0 0 0 28 27 0 0 3
129 106
129 98
121 98
1 1 19 0 0 4224 0 14 29 0 0 2
217 139
228 139
2 0 20 0 0 4096 0 30 0 0 30 2
265 98
273 98
2 1 20 0 0 8320 0 29 18 0 0 4
264 139
273 139
273 98
285 98
1 1 21 0 0 4224 0 15 32 0 0 2
221 86
229 86
1 3 22 0 0 4224 0 17 18 0 0 2
303 73
303 79
1 4 2 0 0 0 0 16 18 0 0 2
303 112
303 105
2 5 23 0 0 8320 0 31 18 0 0 4
321 29
354 29
354 92
321 92
1 0 24 0 0 8320 0 31 0 0 36 3
285 29
273 29
273 86
2 2 24 0 0 0 0 32 18 0 0 2
265 86
285 86
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.05 1e-05 1e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
