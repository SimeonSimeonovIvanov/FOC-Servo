CircuitMaker Text
5.6
Probes: 1
V1_1
Transient Analysis
0 76 60 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 310 10
165 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
333 175 2075 645
9961490 0
0
6 Title:
5 Name:
0
0
0
5
9 I Source~
198 270 60 0 2 5
0 3 2
0
0 0 17264 0
5 250mA
13 0 48 8
3 Is1
20 -10 41 -2
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 1 0 0 0
2 Is
3670 0 0
2
5.8985e-315 0
0
11 Signal Gen~
195 36 64 0 64 64
0 5 4 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1133903872
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 270
20
1 50 0 300 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -300/300V
-32 -30 31 -22
2 V1
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 300 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5616 0 0
2
5.8985e-315 5.32571e-315
0
10 FW Bridge~
219 111 63 0 4 9
0 2 5 3 4
0
0 0 848 90
6 2KBB60
15 -38 57 -30
2 D1
16 -49 30 -41
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 D-37
9

0 1 2 3 4 1 2 3 4 0
88 0 0 256 0 0 0 0
1 D
9323 0 0
2
5.8985e-315 5.30499e-315
0
10 Polar Cap~
219 192 57 0 2 5
0 3 2
0
0 0 848 270
5 100uF
14 4 49 12
2 C1
14 -7 28 1
0
0
11 %D %1 %2 %V
0
0
8 POLAR0.6
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
317 0 0
2
5.8985e-315 5.26354e-315
0
7 Ground~
168 113 126 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
5.8985e-315 0
0
7
2 0 2 0 0 4096 0 4 0 0 5 2
191 64
191 120
1 0 2 0 0 0 0 5 0 0 5 2
113 120
113 120
1 0 3 0 0 8320 0 1 0 0 6 3
270 39
270 4
191 4
2 4 4 0 0 12416 0 2 3 0 0 6
67 69
73 69
73 98
155 98
155 59
145 59
2 1 2 0 0 8320 0 1 3 0 0 4
270 81
270 120
113 120
113 91
3 1 3 0 0 0 0 3 4 0 0 4
113 27
113 4
191 4
191 47
1 2 5 0 0 4224 0 2 3 0 0 2
67 59
81 59
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.1 0.0004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
