CircuitMaker Text
5.6
Probes: 1
R4_2
Transient Analysis
0 346 93 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 130 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
28
10 Capacitor~
219 297 33 0 2 5
0 7 6
0
0 0 848 0
4 10nF
-14 -18 14 -10
2 C1
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
3919 0 0
2
43350.6 27
0
8 Op-Amp5~
219 296 127 0 5 11
0 9 7 14 2 6
0
0 0 848 0
5 AD820
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
9747 0 0
2
43350.6 26
0
11 Signal Gen~
195 30 126 0 64 64
0 11 3 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1127481344 1127481344
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 180 180 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
6 0/360V
-21 -30 21 -22
2 V2
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(180 180 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5310 0 0
2
43350.6 25
0
7 Ground~
168 245 220 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4318 0 0
2
43350.6 24
0
2 +V
167 296 98 0 1 3
0 14
0
0 0 53616 0
4 3.3v
-13 -13 15 -5
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3917 0 0
2
43350.6 23
0
7 Ground~
168 296 150 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7930 0 0
2
43350.6 22
0
11 Signal Gen~
195 31 391 0 64 64
0 16 3 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1073741824 1073741824
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 2 2 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/4V
-15 -30 13 -22
2 V3
-7 -40 7 -32
0
0
36 %D %1 %2 DC 0 SIN(2 2 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6128 0 0
2
43350.6 15
0
7 Ground~
168 298 415 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7346 0 0
2
43350.6 14
0
2 +V
167 298 363 0 1 3
0 19
0
0 0 53616 0
4 3.3v
-13 -13 15 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8577 0 0
2
43350.6 13
0
7 Ground~
168 247 488 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3372 0 0
2
43350.6 12
0
8 Op-Amp5~
219 298 392 0 5 11
0 8 5 19 2 4
0
0 0 848 0
5 AD820
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 256 1 0 0 0
1 U
3741 0 0
2
43350.6 11
0
10 Capacitor~
219 281 182 0 2 5
0 2 9
0
0 0 848 90
4 10nF
12 0 40 8
2 C2
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
5813 0 0
2
43350.6 4
0
10 Capacitor~
219 300 296 0 2 5
0 5 4
0
0 0 848 0
4 10nF
-14 -18 14 -10
2 C3
-7 -28 7 -20
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
3213 0 0
2
43350.6 3
0
10 Capacitor~
219 295 456 0 2 5
0 2 8
0
0 0 848 90
4 10nF
12 0 40 8
2 C4
19 -10 33 -2
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 0 0 0 0
1 C
3694 0 0
2
43350.6 2
0
7 Ground~
168 281 220 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4327 0 0
2
43350.6 1
0
7 Ground~
168 295 488 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8800 0 0
2
43350.6 0
0
11 Resistor:A~
219 297 71 0 2 5
0 7 6
0
0 0 880 0
2 3k
-7 -14 7 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3406 0 0
2
43350.6 21
0
11 Resistor:A~
219 245 184 0 3 5
0 2 9 -1
0
0 0 880 90
2 3k
9 -1 23 7
2 R3
9 -12 23 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6455 0 0
2
43350.6 20
0
11 Resistor:A~
219 216 133 0 2 5
0 12 9
0
0 0 880 0
4 124k
-16 17 12 25
2 R2
-10 7 4 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9319 0 0
2
43350.6 19
0
11 Resistor:A~
219 216 121 0 2 5
0 13 7
0
0 0 880 0
4 124k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3172 0 0
2
43350.6 18
0
11 Resistor:A~
219 146 121 0 2 5
0 3 13
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
38 0 0
2
43350.6 17
0
11 Resistor:A~
219 146 133 0 2 5
0 11 12
0
0 0 880 0
4 224k
-16 17 12 25
2 R7
-10 7 4 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
376 0 0
2
43350.6 16
0
11 Resistor:A~
219 247 457 0 3 5
0 2 8 -1
0
0 0 880 90
4 270k
9 -1 37 7
3 R12
6 -12 27 -4
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6666 0 0
2
43350.6 10
0
11 Resistor:A~
219 299 336 0 2 5
0 5 4
0
0 0 880 0
4 270k
-14 -14 14 -6
3 R13
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9365 0 0
2
43350.6 9
0
11 Resistor:A~
219 147 398 0 2 5
0 16 17
0
0 0 880 0
4 224k
-16 17 12 25
2 R5
-10 7 4 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3251 0 0
2
43350.6 8
0
11 Resistor:A~
219 147 386 0 2 5
0 3 18
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5481 0 0
2
43350.6 7
0
11 Resistor:A~
219 217 386 0 2 5
0 18 5
0
0 0 880 0
4 124k
-14 -14 14 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7788 0 0
2
43350.6 6
0
11 Resistor:A~
219 217 398 0 2 5
0 17 8
0
0 0 880 0
4 124k
-15 18 13 26
3 R10
-13 7 8 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3273 0 0
2
43350.6 5
0
35
0 0 3 0 0 4224 0 0 0 12 27 2
71 131
71 396
2 0 4 0 0 4112 0 13 0 0 30 3
309 296
351 296
351 336
1 0 5 0 0 4112 0 13 0 0 34 3
291 296
247 296
247 336
2 0 6 0 0 4112 0 1 0 0 15 3
306 33
349 33
349 72
1 0 7 0 0 4112 0 1 0 0 16 3
288 33
245 33
245 72
1 1 2 0 0 4112 0 16 14 0 0 2
295 482
295 465
1 1 2 0 0 4240 0 15 12 0 0 2
281 214
281 191
2 0 8 0 0 8336 0 14 0 0 33 3
295 447
295 431
247 431
0 2 9 0 0 4112 0 0 12 17 0 3
245 155
281 155
281 173
0 0 10 0 0 16 0 0 0 0 0 2
150 110
150 110
1 1 11 0 0 12432 0 3 22 0 0 6
61 121
82 121
82 141
106 141
106 133
128 133
2 1 3 0 0 144 0 3 21 0 0 4
61 131
89 131
89 121
128 121
2 1 12 0 0 4240 0 22 19 0 0 2
164 133
198 133
1 2 13 0 0 4240 0 20 21 0 0 2
198 121
164 121
2 5 6 0 0 8336 0 17 2 0 0 4
315 71
349 71
349 127
314 127
0 1 7 0 0 4240 0 0 17 21 0 3
245 121
245 71
279 71
2 0 9 0 0 16 0 18 0 0 20 2
245 166
245 133
1 3 14 0 0 4240 0 5 2 0 0 2
296 107
296 114
1 4 2 0 0 16 0 6 2 0 0 2
296 144
296 140
1 2 9 0 0 4240 0 2 19 0 0 2
278 133
234 133
2 2 7 0 0 16 0 2 20 0 0 2
278 121
234 121
1 1 2 0 0 16 0 4 18 0 0 2
245 214
245 202
2 0 8 0 0 16 0 28 0 0 33 2
235 398
247 398
2 0 5 0 0 16 0 27 0 0 34 2
235 386
247 386
0 0 15 0 0 16 0 0 0 0 0 2
151 375
151 375
1 1 16 0 0 12432 0 7 25 0 0 6
62 386
83 386
83 406
107 406
107 398
129 398
2 1 3 0 0 144 0 7 26 0 0 4
62 396
90 396
90 386
129 386
2 1 17 0 0 4240 0 25 28 0 0 2
165 398
199 398
1 2 18 0 0 4240 0 27 26 0 0 2
199 386
165 386
2 5 4 0 0 8336 0 24 11 0 0 4
317 336
351 336
351 392
316 392
1 3 19 0 0 4240 0 9 11 0 0 2
298 372
298 379
1 4 2 0 0 16 0 8 11 0 0 2
298 409
298 405
2 1 8 0 0 16 0 23 11 0 0 3
247 439
247 398
280 398
1 2 5 0 0 8336 0 24 11 0 0 4
281 336
247 336
247 386
280 386
1 1 2 0 0 16 0 10 23 0 0 2
247 482
247 475
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.1 0.0004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
