CircuitMaker Text
5.6
Probes: 1
Q1_2
Transient Analysis
0 217 97 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 400 10
281 80 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 1
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.823216 0.500000
449 176 2086 949
9961490 0
0
6 Title:
5 Name:
0
0
0
14
11 Signal Gen~
195 36 118 0 64 64
0 5 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1092616192 1075838976 1075419546
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 10 2.5 2.4 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 100m/4.9V
-32 -30 31 -22
2 V3
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(2.5 2.4 10 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
43283.6 9
0
7 Ground~
168 80 171 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6435 0 0
2
43283.6 8
0
2 +V
167 104 32 0 1 3
0 7
0
0 0 53616 0
3 +5V
-11 -14 10 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5283 0 0
2
43283.6 7
0
7 Ground~
168 169 171 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6874 0 0
2
43283.6 6
0
2 +V
167 225 36 0 1 3
0 8
0
0 0 53616 0
3 +5V
-11 -14 10 -6
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5305 0 0
2
43283.6 5
0
2 +V
167 169 77 0 1 3
0 9
0
0 0 53616 0
3 +5V
-11 -14 10 -6
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
34 0 0
2
43283.6 4
0
12 Comparator6~
219 169 107 0 6 13
0 5 3 9 2 6 2
0
0 0 848 0
5 LP311
6 -22 41 -14
2 U1
8 -32 22 -24
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
0
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
88 0 0 0 1 0 0 0
1 U
969 0 0
2
43283.6 3
0
7 Ground~
168 104 171 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8402 0 0
2
43283.6 2
0
12 NPN Trans:B~
219 277 99 0 3 7
0 4 6 2
0
0 0 848 0
8 BC337-16
18 0 74 8
2 Q1
39 -10 53 -2
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 3 2 1 3 2 1 0
81 0 0 0 1 0 0 0
1 Q
3751 0 0
2
43283.6 1
0
7 Ground~
168 282 171 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4292 0 0
2
43283.6 0
0
11 Resistor:A~
219 225 72 0 4 5
0 6 8 0 1
0
0 0 880 90
4 5.1k
7 0 35 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6118 0 0
2
43283.6 13
0
11 Resistor:A~
219 104 140 0 4 5
0 3 2 0 -1
0
0 0 880 270
4 5.1k
8 1 36 9
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
34 0 0
2
43283.6 12
0
11 Resistor:A~
219 104 70 0 3 5
0 7 3 1
0
0 0 880 270
4 5.1k
6 -1 34 7
2 R1
7 -11 21 -3
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6357 0 0
2
43283.6 11
0
11 Resistor:A~
219 282 56 0 2 5
0 3 4
0
0 0 880 270
3 50k
6 0 27 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
319 0 0
2
43283.6 10
0
15
2 0 3 0 0 4096 0 7 0 0 2 2
151 101
104 101
2 1 3 0 0 0 0 13 12 0 0 2
104 88
104 122
1 0 3 0 0 8320 0 14 0 0 1 4
282 38
282 15
145 15
145 101
2 1 4 0 0 4224 0 14 9 0 0 2
282 74
282 81
1 1 5 0 0 4224 0 1 7 0 0 2
67 113
151 113
1 3 2 0 0 4224 0 10 9 0 0 2
282 165
282 117
2 0 6 0 0 4096 0 9 0 0 12 2
259 99
225 99
1 1 7 0 0 4224 0 3 13 0 0 2
104 41
104 52
6 0 2 0 0 0 0 7 0 0 14 4
185 115
196 115
196 143
169 143
2 1 2 0 0 0 0 12 8 0 0 2
104 158
104 165
1 2 8 0 0 4224 0 5 11 0 0 2
225 45
225 54
5 1 6 0 0 4224 0 7 11 0 0 3
185 99
225 99
225 90
1 3 9 0 0 4224 0 6 7 0 0 2
169 86
169 94
1 4 2 0 0 0 0 4 7 0 0 2
169 165
169 120
1 2 2 0 0 0 0 2 1 0 0 3
80 165
80 123
67 123
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.5 0.0002 0.0002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
