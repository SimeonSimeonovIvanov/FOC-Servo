CircuitMaker Text
5.6
Probes: 1
R3_1
Transient Analysis
0 223 86 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 200 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 1
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
12
2 +V
167 111 18 0 1 3
0 5
0
0 0 53616 0
3 +5V
-11 -14 10 -6
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8734 0 0
2
43282.7 11
0
7 Ground~
168 171 157 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7988 0 0
2
43282.7 10
0
7 Ground~
168 80 157 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3217 0 0
2
43282.7 9
0
11 Signal Gen~
195 36 104 0 64 64
0 6 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 1075838976 1075419546
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 1000 2.5 2.4 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 100m/4.9V
-32 -30 31 -22
2 V3
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(2.5 2.4 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3965 0 0
2
43282.7 8
0
2 +V
167 268 19 0 1 3
0 7
0
0 0 53616 0
3 +5V
-11 -14 10 -6
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8239 0 0
2
43282.7 7
0
2 +V
167 171 63 0 1 3
0 8
0
0 0 53616 0
3 +5V
-11 -14 10 -6
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
828 0 0
2
43282.7 6
0
12 Comparator6~
219 171 93 0 6 13
0 6 3 8 2 4 2
0
0 0 848 0
5 LP311
6 -22 41 -14
2 U1
8 -32 22 -24
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
0
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
88 0 0 0 1 0 0 0
1 U
6187 0 0
2
43282.7 5
0
7 Ground~
168 111 157 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7107 0 0
2
43282.7 4
0
11 Resistor:A~
219 220 56 0 2 5
0 3 4
0
0 0 880 270
3 56k
9 0 30 8
2 R4
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6433 0 0
2
43282.7 3
0
11 Resistor:A~
219 268 56 0 4 5
0 4 7 0 1
0
0 0 880 90
4 3.3k
3 0 31 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8559 0 0
2
43282.7 2
0
11 Resistor:A~
219 111 126 0 4 5
0 3 2 0 -1
0
0 0 880 270
2 5k
8 1 22 9
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3674 0 0
2
43282.7 1
0
11 Resistor:A~
219 111 56 0 3 5
0 5 3 1
0
0 0 880 270
2 5k
9 0 23 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5697 0 0
2
43282.7 0
0
13
1 0 3 0 0 8336 0 9 0 0 4 4
220 38
220 26
141 26
141 87
2 0 4 0 0 4112 0 9 0 0 11 2
220 74
220 85
1 1 5 0 0 4240 0 1 12 0 0 2
111 27
111 38
2 0 3 0 0 16 0 7 0 0 5 2
153 87
111 87
2 1 3 0 0 16 0 12 11 0 0 2
111 74
111 108
1 1 6 0 0 4240 0 4 7 0 0 2
67 99
153 99
6 0 2 0 0 12304 0 7 0 0 13 4
187 101
211 101
211 129
171 129
1 2 2 0 0 4112 0 3 4 0 0 3
80 151
80 109
67 109
2 1 2 0 0 16 0 11 8 0 0 2
111 144
111 151
1 2 7 0 0 4240 0 5 10 0 0 2
268 28
268 38
5 1 4 0 0 4240 0 7 10 0 0 3
187 85
268 85
268 74
1 3 8 0 0 4240 0 6 7 0 0 2
171 72
171 80
1 4 2 0 0 4240 0 2 7 0 0 2
171 151
171 106
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
