CircuitMaker Text
5.6
Probes: 1
U1_1
Transient Analysis
0 117 126 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 210 10
176 79 1918 521
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 1
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.520213 0.500000
344 175 2086 664
9961490 0
0
6 Title:
5 Name:
0
0
0
16
7 Ground~
168 333 57 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
363 0 0
2
43315 10
0
7 Ground~
168 108 187 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8132 0 0
2
43315 9
0
12 Comparator6~
219 182 80 0 6 13
0 9 8 11 7 5 7
0
0 0 848 0
5 LP311
6 -22 41 -14
2 U1
8 -32 22 -24
0
0
23 %D %1 %2 %3 %4 %5 %6 %S
0
0
0
13

0 1 2 3 4 5 6 1 2 3
4 5 6 0
88 0 0 0 1 0 0 0
1 U
65 0 0
2
43315 8
0
2 +V
167 182 122 0 1 3
0 7
0
0 0 53616 180
4 -15V
-13 -1 15 7
2 V1
10 -12 24 -4
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6609 0 0
2
43315 7
0
2 +V
167 182 50 0 1 3
0 11
0
0 0 53616 0
4 +15V
-14 -14 14 -6
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8995 0 0
2
43315 6
0
2 +V
167 248 16 0 1 3
0 10
0
0 0 53616 0
4 +15V
-14 -13 14 -5
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3918 0 0
2
43315 5
0
11 Signal Gen~
195 28 79 0 64 64
0 8 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1120403456 0 1092616192
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 100 0 10 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -10/10V
-25 -30 24 -22
2 V3
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 10 100 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
7519 0 0
2
43315 4
0
7 Ground~
168 72 110 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
377 0 0
2
43315 3
0
14 Opto Isolator~
173 379 60 0 4 9
0 2 6 3 4
0
0 0 880 0
6 OP4N25
-21 -28 21 -20
2 U2
-7 -38 7 -30
0
0
17 %D %1 %2 %3 %4 %S
0
0
4 DIP6
9

0 1 2 5 4 1 2 5 4 0
88 0 0 0 1 0 0 0
1 U
8816 0 0
2
43315 2
0
7 Ground~
168 417 131 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -28 14 -20
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3877 0 0
2
43315 1
0
2 +V
167 417 32 0 1 3
0 3
0
0 0 53616 0
5 +3.3V
-17 -14 18 -6
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
926 0 0
2
43315 0
0
11 Resistor:A~
219 296 72 0 2 5
0 6 5
0
0 0 880 180
3 10k
-10 -14 11 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7262 0 0
2
43315 15
0
11 Resistor:A~
219 108 100 0 2 5
0 5 9
0
0 0 880 270
3 20k
8 0 29 8
2 R1
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5267 0 0
2
43315 14
0
11 Resistor:A~
219 108 156 0 4 5
0 9 2 0 -1
0
0 0 880 270
3 120
9 0 30 8
2 R2
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8838 0 0
2
43315 13
0
11 Resistor:A~
219 248 47 0 4 5
0 5 10 0 1
0
0 0 880 90
3 10k
6 0 27 8
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7159 0 0
2
43315 12
0
11 Resistor:A~
219 417 100 0 4 5
0 4 2 0 -1
0
0 0 880 270
4 3.3k
6 0 34 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5812 0 0
2
43315 11
0
17
1 3 3 0 0 8336 0 11 9 0 0 3
417 41
417 48
405 48
1 2 2 0 0 4112 0 10 16 0 0 2
417 125
417 118
1 4 4 0 0 8336 0 16 9 0 0 3
417 82
417 72
405 72
1 1 2 0 0 8208 0 1 9 0 0 3
333 51
333 48
351 48
2 0 5 0 0 4112 0 12 0 0 15 2
278 72
223 72
1 0 5 0 0 16 0 15 0 0 5 2
248 65
248 72
2 1 6 0 0 4240 0 9 12 0 0 2
351 72
314 72
6 0 7 0 0 12432 0 3 0 0 17 4
198 88
222 88
222 102
182 102
1 2 8 0 0 4240 0 7 3 0 0 2
59 74
164 74
1 2 2 0 0 4240 0 8 7 0 0 3
72 104
72 84
59 84
2 1 2 0 0 16 0 14 2 0 0 2
108 174
108 181
1 0 9 0 0 12432 0 3 0 0 13 4
164 86
149 86
149 126
108 126
2 1 9 0 0 16 0 13 14 0 0 2
108 118
108 138
1 2 10 0 0 4240 0 6 15 0 0 2
248 25
248 29
5 1 5 0 0 12432 0 3 13 0 0 5
198 72
223 72
223 12
108 12
108 82
1 3 11 0 0 4240 0 5 3 0 0 2
182 59
182 67
1 4 7 0 0 16 0 4 3 0 0 2
182 107
182 93
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.05 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
