CircuitMaker Text
5.6
Probes: 1
U1B_7
Transient Analysis
0 685 88 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 79 1918 540
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 2 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
30
11 Signal Gen~
195 399 112 0 64 64
0 15 16 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846080 1075838976 1065353216
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 44315892
20
0 1000 2.5 1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
8 1.5/3.5V
-29 -30 27 -22
2 V4
-8 -40 6 -32
0
0
31 %D %1 %2 DC 0 SIN(2.5 1 1k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3409 0 0
2
5.89888e-315 0
0
11 Signal Gen~
195 43 290 0 64 64
0 3 4 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846080 1075838976 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 34
20
0 1000 2.5 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 2/3V
-15 -30 13 -22
2 V7
-8 -40 6 -32
0
0
34 %D %1 %2 DC 0 SIN(2.5 500m 1k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3951 0 0
2
5.89888e-315 0
0
8 Op-Amp5~
219 284 289 0 5 11
0 6 7 8 2 9
0
0 0 848 0
5 LM358
11 6 46 14
3 U2A
12 -13 33 -5
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 2 0
1 U
8885 0 0
2
5.89888e-315 5.34643e-315
0
2 +V
167 237 363 0 1 3
0 5
0
0 0 54128 180
4 1.65
-12 12 16 20
5 Vref3
-15 1 20 9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3780 0 0
2
5.89888e-315 5.32571e-315
0
7 Ground~
168 284 315 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9265 0 0
2
5.89888e-315 5.26354e-315
0
2 +V
167 284 256 0 1 3
0 8
0
0 0 54128 0
2 10
-6 -13 8 -5
2 V6
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9442 0 0
2
5.89888e-315 0
0
2 +V
167 638 145 0 1 3
0 12
0
0 0 54128 180
3 -10
-8 1 13 9
2 V5
-3 11 11 19
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9424 0 0
2
43599 0
0
8 Op-Amp5~
219 638 111 0 5 11
0 18 19 20 12 21
0
0 0 848 0
5 LM358
11 6 46 14
3 U1B
12 -13 33 -5
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
9968 0 0
2
5.89888e-315 0
0
2 +V
167 591 185 0 1 3
0 17
0
0 0 54128 180
2 0v
-4 12 10 20
5 Vref2
-15 1 20 9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
9281 0 0
2
5.89888e-315 5.26354e-315
0
2 +V
167 638 78 0 1 3
0 20
0
0 0 54128 0
2 10
-6 -13 8 -5
2 V3
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8464 0 0
2
5.89888e-315 5.32571e-315
0
2 +V
167 287 69 0 1 3
0 25
0
0 0 54128 0
2 10
-6 -13 8 -5
2 V2
-7 -23 7 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7168 0 0
2
5.89888e-315 5.34643e-315
0
7 Ground~
168 287 128 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3171 0 0
2
5.89888e-315 5.3568e-315
0
11 Signal Gen~
195 48 103 0 64 64
0 13 14 2 86 -10 10 0 0 0
0 0 0 0 0 0 0 1148846080 0 1056964608
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
0 1000 0 0.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -500m/500mV
-39 -30 38 -22
2 V1
-8 -40 6 -32
0
0
32 %D %1 %2 DC 0 SIN(0 500m 1k 0 0)
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
5.89888e-315 5.36716e-315
0
2 +V
167 240 176 0 1 3
0 22
0
0 0 54128 180
4 1.65
-12 12 16 20
5 Vref1
-15 1 20 9
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6435 0 0
2
5.89888e-315 5.37752e-315
0
8 Op-Amp5~
219 287 102 0 5 11
0 23 24 25 2 26
0
0 0 848 0
5 LM358
11 6 46 14
3 U1A
12 -13 33 -5
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
5283 0 0
2
5.89888e-315 5.38788e-315
0
11 Resistor:A~
219 146 290 0 2 5
0 3 4
0
0 0 880 90
3 120
7 0 28 8
3 R15
8 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6874 0 0
2
5.89888e-315 5.39306e-315
0
11 Resistor:A~
219 198 295 0 2 5
0 3 6
0
0 0 880 0
2 3k
-6 16 8 24
3 R14
-14 6 7 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5305 0 0
2
5.89888e-315 5.38788e-315
0
11 Resistor:A~
219 237 325 0 3 5
0 5 6 1
0
0 0 880 90
2 3k
10 0 24 8
3 R13
8 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
34 0 0
2
5.89888e-315 5.37752e-315
0
11 Resistor:A~
219 198 283 0 2 5
0 4 7
0
0 0 880 0
2 3k
-6 -14 8 -6
3 R12
-9 -24 12 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
969 0 0
2
5.89888e-315 5.36716e-315
0
11 Resistor:A~
219 281 219 0 2 5
0 7 9
0
0 0 880 0
2 3k
-6 -14 8 -6
3 R11
-9 -24 12 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8402 0 0
2
5.89888e-315 5.3568e-315
0
11 Resistor:A~
219 500 112 0 2 5
0 15 16
0
0 0 880 90
3 120
7 0 28 8
3 R10
8 -10 29 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3751 0 0
2
5.89888e-315 5.39306e-315
0
11 Resistor:A~
219 552 117 0 2 5
0 15 18
0
0 0 880 0
2 3k
-6 16 8 24
2 R9
-11 6 3 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4292 0 0
2
5.89888e-315 5.39824e-315
0
11 Resistor:A~
219 591 147 0 3 5
0 17 18 1
0
0 0 880 90
4 1.5k
3 0 31 8
2 R8
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6118 0 0
2
5.89888e-315 5.40342e-315
0
11 Resistor:A~
219 552 105 0 2 5
0 16 19
0
0 0 880 0
2 3k
-6 -14 8 -6
2 R5
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
34 0 0
2
5.89888e-315 5.4086e-315
0
11 Resistor:A~
219 635 41 0 2 5
0 19 21
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R4
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6357 0 0
2
5.89888e-315 5.41378e-315
0
11 Resistor:A~
219 284 32 0 2 5
0 24 26
0
0 0 880 0
2 3k
-6 -14 8 -6
2 R7
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
319 0 0
2
5.89888e-315 5.41896e-315
0
11 Resistor:A~
219 201 96 0 2 5
0 14 24
0
0 0 880 0
4 1.5k
-13 -14 15 -6
2 R6
-6 -24 8 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3976 0 0
2
5.89888e-315 5.42414e-315
0
11 Resistor:A~
219 240 138 0 3 5
0 22 23 1
0
0 0 880 90
2 3k
10 0 24 8
2 R1
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7634 0 0
2
5.89888e-315 5.42933e-315
0
11 Resistor:A~
219 201 108 0 2 5
0 13 23
0
0 0 880 0
4 1.5k
-13 16 15 24
2 R2
-11 6 3 14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
523 0 0
2
5.89888e-315 5.43192e-315
0
11 Resistor:A~
219 149 103 0 2 5
0 13 14
0
0 0 880 90
3 120
7 0 28 8
2 R3
11 -10 25 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6748 0 0
2
5.89888e-315 5.43451e-315
0
38
1 0 3 0 0 12416 0 2 0 0 5 4
74 285
94 285
94 313
147 313
2 0 4 0 0 12416 0 2 0 0 4 4
74 295
108 295
108 265
146 265
1 1 5 0 0 4224 0 4 18 0 0 2
237 348
237 343
2 1 4 0 0 0 0 16 19 0 0 5
146 272
146 265
174 265
174 283
180 283
1 1 3 0 0 0 0 17 16 0 0 5
180 295
174 295
174 313
146 313
146 308
2 0 6 0 0 4096 0 18 0 0 7 2
237 307
237 295
2 1 6 0 0 4224 0 17 3 0 0 2
216 295
266 295
1 4 2 0 0 4224 0 5 3 0 0 2
284 309
284 302
1 0 7 0 0 8320 0 20 0 0 10 3
263 219
237 219
237 283
2 2 7 0 0 0 0 19 3 0 0 2
216 283
266 283
1 3 8 0 0 4224 0 6 3 0 0 2
284 265
284 276
5 2 9 0 0 8320 0 3 20 0 0 4
302 289
329 289
329 219
299 219
0 0 10 0 0 0 0 0 0 0 0 2
448 160
448 160
0 0 11 0 0 4224 0 0 0 0 0 2
500 135
448 135
1 4 12 0 0 4224 0 7 8 0 0 2
638 130
638 124
1 0 13 0 0 12416 0 13 0 0 31 4
79 98
97 98
97 126
150 126
2 0 14 0 0 12416 0 13 0 0 30 4
79 108
111 108
111 78
149 78
1 0 15 0 0 12416 0 1 0 0 22 4
430 107
448 107
448 135
500 135
2 0 16 0 0 12416 0 1 0 0 21 4
430 117
463 117
463 87
500 87
1 1 17 0 0 4224 0 9 23 0 0 2
591 170
591 165
2 1 16 0 0 0 0 21 24 0 0 5
500 94
500 87
528 87
528 105
534 105
1 1 15 0 0 0 0 22 21 0 0 5
534 117
528 117
528 135
500 135
500 130
2 0 18 0 0 4096 0 23 0 0 24 2
591 129
591 117
2 1 18 0 0 4224 0 22 8 0 0 2
570 117
620 117
1 0 19 0 0 8320 0 25 0 0 26 3
617 41
591 41
591 105
2 2 19 0 0 0 0 24 8 0 0 2
570 105
620 105
1 3 20 0 0 4224 0 10 8 0 0 2
638 87
638 98
5 2 21 0 0 8320 0 8 25 0 0 4
656 111
683 111
683 41
653 41
1 1 22 0 0 4224 0 14 28 0 0 2
240 161
240 156
2 1 14 0 0 0 0 30 27 0 0 5
149 85
149 78
177 78
177 96
183 96
1 1 13 0 0 0 0 29 30 0 0 5
183 108
177 108
177 126
149 126
149 121
2 0 23 0 0 4096 0 28 0 0 33 2
240 120
240 108
2 1 23 0 0 4224 0 29 15 0 0 2
219 108
269 108
1 4 2 0 0 0 0 12 15 0 0 2
287 122
287 115
1 0 24 0 0 8320 0 26 0 0 36 3
266 32
240 32
240 96
2 2 24 0 0 0 0 27 15 0 0 2
219 96
269 96
1 3 25 0 0 4224 0 11 15 0 0 2
287 78
287 89
5 2 26 0 0 8320 0 15 26 0 0 4
305 102
332 102
332 32
302 32
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
