CircuitMaker Text
5.6
Probes: 10
r2[p]
AC Analysis
0 117 130 65280
r2[p]
DC Sweep
0 117 130 65280
r2[p]
Operating Point
0 117 130 65280
r2[p]
Transient Analysis
0 117 130 65280
r2[p]
Fourier Analysis
0 117 130 65280
r21[p]
AC Analysis
1 115 319 65535
r21[p]
DC Sweep
1 115 319 65535
r21[p]
Operating Point
1 115 319 65535
r21[p]
Transient Analysis
1 115 319 65535
r21[p]
Fourier Analysis
1 115 319 65535
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 120 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
50
10 Op-Amp5:A~
219 331 96 0 5 11
0 28 27 34 2 33
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
754 0 0
2
43282.7 21
0
7 Ground~
168 331 120 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9767 0 0
2
43282.7 20
0
2 +V
167 331 44 0 1 3
0 34
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
7978 0 0
2
43282.7 19
0
7 Ground~
168 284 24 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3142 0 0
2
43282.7 18
0
11 Signal Gen~
195 41 107 0 64 64
0 32 31 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1133903872 1133903872
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 300 300 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
6 0/600V
-22 -30 20 -22
2 V2
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(300 300 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3284 0 0
2
43282.7 17
0
5 SAVE-
218 117 130 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
659 0 0
2
43282.7 16
0
5 SAVE-
218 115 319 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
3800 0 0
2
43282.7 15
0
11 Signal Gen~
195 39 296 0 64 64
0 24 23 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1127481344 1127481344
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 180 180 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
6 0/360V
-22 -30 20 -22
2 V7
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(180 180 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
6792 0 0
2
43282.7 14
0
7 Ground~
168 282 213 0 1 3
0 2
0
0 0 53360 180
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3701 0 0
2
43282.7 13
0
2 +V
167 329 233 0 1 3
0 26
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6316 0 0
2
43282.7 12
0
7 Ground~
168 329 309 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8734 0 0
2
43282.7 11
0
10 Op-Amp5:A~
219 329 285 0 5 11
0 20 19 26 2 25
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U4
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
7988 0 0
2
43282.7 10
0
11 Signal Gen~
195 457 111 0 64 64
0 18 17 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1075838976 1075838976
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 2.5 2.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/5V
-15 -30 13 -22
2 V5
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(2.5 2.5 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3217 0 0
2
43282.7 9
0
7 Ground~
168 688 22 0 1 3
0 2
0
0 0 53360 180
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3965 0 0
2
43282.7 8
0
2 +V
167 735 52 0 1 3
0 15
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8239 0 0
2
43282.7 7
0
7 Ground~
168 735 118 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
828 0 0
2
43282.7 6
0
10 Op-Amp5:A~
219 735 93 0 5 11
0 14 12 15 2 13
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U3
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
6187 0 0
2
43282.7 5
0
10 Op-Amp5:A~
219 723 283 0 5 11
0 6 4 7 2 5
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 1 0 0 0
1 U
7107 0 0
2
43282.7 4
0
7 Ground~
168 723 308 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6433 0 0
2
43282.7 3
0
2 +V
167 723 242 0 1 3
0 7
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
8559 0 0
2
43282.7 2
0
7 Ground~
168 676 212 0 1 3
0 2
0
0 0 53360 180
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3674 0 0
2
43282.7 1
0
11 Signal Gen~
195 445 301 0 64 64
0 10 9 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1142292480
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 26
20
1 50 0 600 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -600/600V
-32 -30 31 -22
2 V4
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 600 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
5697 0 0
2
43282.7 0
0
11 Resistor:A~
219 284 59 0 3 5
0 2 28 -1
0
0 0 880 270
4 6.8k
7 1 35 9
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3805 0 0
2
43282.7 49
0
11 Resistor:A~
219 330 163 0 2 5
0 33 27
0
0 0 880 180
4 6.8k
-16 -14 12 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5219 0 0
2
43282.7 48
0
11 Resistor:A~
219 155 107 0 2 5
0 30 29
0
0 0 880 90
3 56k
8 0 29 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3795 0 0
2
43282.7 47
0
11 Resistor:A~
219 117 130 0 2 5
0 31 30
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3637 0 0
2
43282.7 46
0
11 Resistor:A~
219 118 83 0 2 5
0 32 29
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3226 0 0
2
43282.7 45
0
11 Resistor:A~
219 201 85 0 2 5
0 29 28
0
0 0 880 0
4 124k
-14 -14 14 -6
3 R16
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6966 0 0
2
43282.7 44
0
11 Resistor:A~
219 198 128 0 2 5
0 30 27
0
0 0 880 0
4 124k
-14 -14 14 -6
3 R17
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9796 0 0
2
43282.7 43
0
11 Resistor:A~
219 196 317 0 2 5
0 22 19
0
0 0 880 0
4 124k
-14 -14 14 -6
3 R18
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5952 0 0
2
43282.7 42
0
11 Resistor:A~
219 199 274 0 2 5
0 21 20
0
0 0 880 0
4 124k
-14 -14 14 -6
3 R19
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3649 0 0
2
43282.7 41
0
11 Resistor:A~
219 116 272 0 2 5
0 24 21
0
0 0 880 0
4 224k
-14 -14 14 -6
3 R20
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3716 0 0
2
43282.7 40
0
11 Resistor:A~
219 115 319 0 2 5
0 23 22
0
0 0 880 0
4 224k
-14 -14 14 -6
3 R21
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4797 0 0
2
43282.7 39
0
11 Resistor:A~
219 153 296 0 2 5
0 22 21
0
0 0 880 90
3 56k
8 0 29 8
3 R22
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4681 0 0
2
43282.7 38
0
11 Resistor:A~
219 328 352 0 2 5
0 25 19
0
0 0 880 180
3 11k
-13 -14 8 -6
3 R23
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9730 0 0
2
43282.7 37
0
11 Resistor:A~
219 282 248 0 3 5
0 2 20 -1
0
0 0 880 270
3 11k
10 1 31 9
3 R24
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9874 0 0
2
43282.7 36
0
11 Resistor:A~
219 734 161 0 2 5
0 13 12
0
0 0 880 180
4 200k
-14 -14 14 -6
3 R15
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
364 0 0
2
43282.7 35
0
11 Resistor:A~
219 688 57 0 3 5
0 2 14 -1
0
0 0 880 270
4 200k
9 1 37 9
3 R14
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3656 0 0
2
43282.7 34
0
11 Resistor:A~
219 629 87 0 2 5
0 16 14
0
0 0 880 0
4 10k2
-13 -14 15 -6
3 R26
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3131 0 0
2
43282.7 33
0
11 Resistor:A~
219 627 134 0 2 5
0 11 12
0
0 0 880 0
4 10k2
-13 -14 15 -6
3 R25
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6772 0 0
2
43282.7 32
0
11 Resistor:A~
219 536 134 0 2 5
0 17 11
0
0 0 880 0
4 224k
-14 -14 14 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9557 0 0
2
43282.7 31
0
11 Resistor:A~
219 537 87 0 2 5
0 18 16
0
0 0 880 0
4 224k
-14 -14 14 -6
3 R11
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
5789 0 0
2
43282.7 30
0
11 Resistor:A~
219 525 277 0 2 5
0 10 8
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7328 0 0
2
43282.7 29
0
11 Resistor:A~
219 524 324 0 2 5
0 9 3
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4799 0 0
2
43282.7 28
0
11 Resistor:A~
219 615 324 0 2 5
0 3 4
0
0 0 880 0
4 10k2
-14 -14 14 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9196 0 0
2
43282.7 27
0
11 Resistor:A~
219 617 277 0 2 5
0 8 6
0
0 0 880 0
4 10k2
-14 -14 14 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3857 0 0
2
43282.7 26
0
11 Resistor:A~
219 676 247 0 3 5
0 2 6 -1
0
0 0 880 270
4 200k
9 1 37 9
3 R10
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7125 0 0
2
43282.7 25
0
11 Resistor:A~
219 722 351 0 2 5
0 5 4
0
0 0 880 180
4 200k
-14 -14 14 -6
3 R27
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3641 0 0
2
43282.7 24
0
11 Resistor:A~
219 562 302 0 2 5
0 3 8
0
0 0 880 90
3 56k
8 0 29 8
3 R28
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9821 0 0
2
43282.7 23
0
11 Resistor:A~
219 574 110 0 2 5
0 11 16
0
0 0 880 90
3 56k
8 0 29 8
3 R13
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3187 0 0
2
43282.7 22
0
56
1 0 3 0 0 4240 0 45 0 0 12 2
597 324
561 324
2 0 4 0 0 4112 0 45 0 0 4 2
633 324
676 324
5 1 5 0 0 8336 0 18 48 0 0 4
741 283
756 283
756 351
740 351
2 2 4 0 0 8336 0 48 18 0 0 4
704 351
676 351
676 289
705 289
1 1 2 0 0 4240 0 21 47 0 0 2
676 220
676 229
2 0 6 0 0 4240 0 46 0 0 7 2
635 277
676 277
1 2 6 0 0 16 0 18 47 0 0 5
705 277
676 277
676 278
676 278
676 265
1 3 7 0 0 4240 0 20 18 0 0 2
723 251
723 270
1 4 2 0 0 16 0 19 18 0 0 2
723 302
723 296
1 0 8 0 0 4240 0 46 0 0 11 2
599 277
562 277
2 2 8 0 0 16 0 43 49 0 0 3
543 277
562 277
562 284
2 1 3 0 0 16 0 44 49 0 0 3
542 324
562 324
562 320
1 2 9 0 0 8336 0 44 22 0 0 4
506 324
491 324
491 306
476 306
1 1 10 0 0 8336 0 22 43 0 0 4
476 296
491 296
491 277
507 277
1 0 11 0 0 4240 0 40 0 0 26 2
609 134
573 134
2 0 12 0 0 4112 0 40 0 0 18 2
645 134
688 134
5 1 13 0 0 8336 0 17 37 0 0 4
753 93
768 93
768 161
752 161
2 2 12 0 0 8336 0 37 17 0 0 4
716 161
688 161
688 99
717 99
1 1 2 0 0 16 0 14 38 0 0 2
688 30
688 39
2 0 14 0 0 4240 0 39 0 0 21 2
647 87
688 87
1 2 14 0 0 16 0 17 38 0 0 5
717 87
688 87
688 88
688 88
688 75
1 3 15 0 0 4240 0 15 17 0 0 2
735 61
735 80
1 4 2 0 0 16 0 16 17 0 0 2
735 112
735 106
1 0 16 0 0 4240 0 39 0 0 25 2
611 87
574 87
2 2 16 0 0 16 0 42 50 0 0 3
555 87
574 87
574 92
2 1 11 0 0 16 0 41 50 0 0 3
554 134
574 134
574 128
1 2 17 0 0 8336 0 41 13 0 0 4
518 134
503 134
503 116
488 116
1 1 18 0 0 8336 0 13 42 0 0 4
488 106
503 106
503 87
519 87
2 0 19 0 0 4240 0 30 0 0 38 2
214 317
282 317
2 0 20 0 0 4240 0 31 0 0 40 2
217 274
282 274
1 0 21 0 0 8336 0 31 0 0 33 3
181 274
181 272
153 272
1 0 22 0 0 8336 0 30 0 0 34 3
178 317
178 319
153 319
2 2 21 0 0 16 0 32 34 0 0 3
134 272
153 272
153 278
2 1 22 0 0 16 0 33 34 0 0 3
133 319
153 319
153 314
1 2 23 0 0 8336 0 33 8 0 0 4
97 319
82 319
82 301
70 301
1 1 24 0 0 8336 0 8 32 0 0 4
70 291
82 291
82 272
98 272
5 1 25 0 0 8336 0 12 35 0 0 4
347 285
362 285
362 352
346 352
2 2 19 0 0 16 0 35 12 0 0 4
310 352
282 352
282 291
311 291
1 1 2 0 0 16 0 9 36 0 0 2
282 221
282 230
1 2 20 0 0 16 0 12 36 0 0 3
311 279
282 279
282 266
1 3 26 0 0 4240 0 10 12 0 0 2
329 242
329 272
1 4 2 0 0 16 0 11 12 0 0 2
329 303
329 298
2 0 27 0 0 4240 0 29 0 0 52 2
216 128
284 128
2 0 28 0 0 4240 0 28 0 0 54 2
219 85
284 85
1 0 29 0 0 8336 0 28 0 0 47 3
183 85
183 83
155 83
1 0 30 0 0 8336 0 29 0 0 48 3
180 128
180 130
155 130
2 2 29 0 0 16 0 27 25 0 0 3
136 83
155 83
155 89
2 1 30 0 0 16 0 26 25 0 0 3
135 130
155 130
155 125
1 2 31 0 0 8336 0 26 5 0 0 4
99 130
84 130
84 112
72 112
1 1 32 0 0 8336 0 5 27 0 0 4
72 102
84 102
84 83
100 83
5 1 33 0 0 8336 0 1 24 0 0 4
349 96
364 96
364 163
348 163
2 2 27 0 0 16 0 24 1 0 0 4
312 163
284 163
284 102
313 102
1 1 2 0 0 16 0 4 23 0 0 2
284 32
284 41
1 2 28 0 0 16 0 1 23 0 0 3
313 90
284 90
284 77
1 3 34 0 0 4240 0 3 1 0 0 2
331 53
331 83
1 4 2 0 0 16 0 2 1 0 0 2
331 114
331 109
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.1 0.0004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
