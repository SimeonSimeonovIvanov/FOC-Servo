CircuitMaker Text
5.6
Probes: 5
U1B_7
AC Analysis
1 294 89 65535
U1B_7
DC Sweep
1 294 89 65535
U1B_7
Operating Point
1 294 89 65535
U1B_7
Fourier Analysis
1 294 89 65535
U1B_7
Transient Analysis
0 275 90 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 230 10
176 83 1918 1019
8  5.000 V
8  5.000 V
3 GND
0 0
24 100 0 2 1
20 Package,Description,
28 C:\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 179 2086 647
9961490 0
0
6 Title:
5 Name:
0
0
0
15
5 SAVE-
218 293 86 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
6901 0 0
2
42769 8
0
2 +V
167 127 29 0 1 3
0 6
0
0 0 53616 0
4 3.3V
-13 -14 15 -6
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
842 0 0
2
42769 7
0
2 +V
167 235 64 0 1 3
0 10
0
0 0 53616 0
4 3.3V
-13 -14 15 -6
2 V5
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3277 0 0
2
42769 6
0
8 Op-Amp5~
219 235 91 0 5 11
0 7 9 10 2 8
0
0 0 848 0
6 OP284E
12 -25 54 -17
3 U1B
22 -35 43 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
4212 0 0
2
42769 5
0
7 Ground~
168 235 117 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4720 0 0
2
42769 4
0
2 +V
167 144 87 0 1 3
0 5
0
0 0 53616 90
4 1.8V
-12 -16 16 -8
2 V7
-6 -28 8 -20
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5551 0 0
2
42769 3
0
7 Ground~
168 265 179 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6986 0 0
2
42769 2
0
11 Signal Gen~
195 31 130 0 64 64
0 3 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1092616192 0 1092616192
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 10 0 10 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 -10/10V
-23 -30 26 -22
2 V6
-7 -40 7 -32
0
0
37 %D %1 %2 DC 0 SIN(0 10 10 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
8745 0 0
2
42769 1
0
7 Ground~
168 79 154 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9592 0 0
2
42769 0
0
11 Resistor:A~
219 174 97 0 3 5
0 6 7 1
0
0 0 880 0
3 51k
-12 14 9 22
2 R4
-12 5 2 13
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
8748 0 0
2
42769 14
0
11 Resistor:A~
219 174 85 0 3 5
0 5 9 1
0
0 0 880 0
3 51k
-10 -14 11 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7168 0 0
2
42769 13
0
11 Resistor:A~
219 234 28 0 2 5
0 9 8
0
0 0 880 0
3 51k
-10 -14 11 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
631 0 0
2
42769 12
0
11 Resistor:A~
219 206 138 0 2 5
0 4 7
0
0 0 880 90
3 51k
-29 1 -8 9
2 R8
-28 -10 -14 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
9466 0 0
2
42769 11
0
11 Resistor:A~
219 160 168 0 2 5
0 4 3
0
0 0 880 180
4 6.2k
-15 -14 13 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3266 0 0
2
42769 10
0
11 Resistor:A~
219 236 168 0 3 5
0 2 4 -1
0
0 0 880 180
4 1.1k
-14 -14 14 -6
3 R10
-11 -24 10 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7693 0 0
2
42769 9
0
14
1 2 3 0 0 4240 0 8 14 0 0 4
62 125
127 125
127 168
142 168
2 1 2 0 0 4240 0 8 9 0 0 3
62 135
79 135
79 148
1 1 2 0 0 16 0 15 7 0 0 3
254 168
265 168
265 173
1 0 4 0 0 4240 0 14 0 0 5 2
178 168
206 168
2 1 4 0 0 16 0 15 13 0 0 3
218 168
206 168
206 156
1 1 5 0 0 4240 0 6 11 0 0 2
155 85
156 85
1 1 6 0 0 8336 0 10 2 0 0 3
156 97
127 97
127 38
2 0 7 0 0 4112 0 13 0 0 12 2
206 120
206 97
2 5 8 0 0 8336 0 12 4 0 0 4
252 28
294 28
294 91
253 91
1 0 9 0 0 8336 0 12 0 0 11 3
216 28
206 28
206 85
2 2 9 0 0 16 0 11 4 0 0 2
192 85
217 85
2 1 7 0 0 4240 0 10 4 0 0 2
192 97
217 97
1 4 2 0 0 16 0 5 4 0 0 2
235 111
235 104
1 3 10 0 0 4240 0 3 4 0 0 2
235 73
235 78
0
0
2065 2 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1 0.002 0.002
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
