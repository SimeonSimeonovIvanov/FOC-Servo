CircuitMaker Text
5.6
Probes: 1
R27_1
Transient Analysis
0 1041 602 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
300 290 30 120 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 2086 645
9961490 0
0
6 Title:
5 Name:
0
0
0
50
11 Signal Gen~
195 733 582 0 64 64
0 10 9 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 0 1142292480
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 50 0 600 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
9 -600/600V
-32 -30 31 -22
2 V4
-7 -40 7 -32
0
0
38 %D %1 %2 DC 0 SIN(0 600 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
7542 0 0
2
43274.8 11
0
7 Ground~
168 964 493 0 1 3
0 2
0
0 0 53360 180
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9283 0 0
2
43274.8 10
0
2 +V
167 1011 523 0 1 3
0 7
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V3
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3600 0 0
2
43274.8 9
0
7 Ground~
168 1011 589 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
8274 0 0
2
43274.8 8
0
10 Op-Amp5:A~
219 1011 564 0 5 11
0 6 4 7 2 5
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U2
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 0 0 0 0
1 U
3329 0 0
2
43274.8 7
0
10 Op-Amp5:A~
219 1023 374 0 5 11
0 14 12 15 2 13
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U3
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 0 0 0 0
1 U
3509 0 0
2
43274.8 4
0
7 Ground~
168 1023 399 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
90 0 0
2
43274.8 3
0
2 +V
167 1023 333 0 1 3
0 15
0
0 0 54256 0
2 5V
-8 -22 6 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
5259 0 0
2
43274.8 2
0
7 Ground~
168 976 303 0 1 3
0 2
0
0 0 53360 180
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6548 0 0
2
43274.8 1
0
11 Signal Gen~
195 745 392 0 64 64
0 18 17 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1075838976 1075838976
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 6721428
20
1 50 2.5 2.5 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
4 0/5V
-15 -30 13 -22
2 V5
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(2.5 2.5 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9326 0 0
2
43274.8 0
0
10 Op-Amp5:A~
219 617 566 0 5 11
0 20 19 26 2 25
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U4
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 0 0 0 0
1 U
5634 0 0
2
43274.8 5
0
7 Ground~
168 617 590 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7902 0 0
2
43274.8 4
0
2 +V
167 617 514 0 1 3
0 26
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V8
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
6805 0 0
2
43274.8 3
0
7 Ground~
168 570 494 0 1 3
0 2
0
0 0 53360 180
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6198 0 0
2
43274.8 2
0
11 Signal Gen~
195 327 577 0 64 64
0 24 23 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1127481344 1127481344
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 18
20
1 50 180 180 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
6 0/360V
-22 -30 20 -22
2 V7
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(180 180 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
9216 0 0
2
43274.8 1
0
5 SAVE-
218 403 600 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 B
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
4 SAVE
9719 0 0
2
43274.8 0
0
5 SAVE-
218 405 411 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57552 0
1 A
3 -26 10 -18
0
0
0
0
0
0
0
3

0 0 0 0
0 0 0 0 0 0 0 0
4 SAVE
3781 0 0
2
43274.8 0
0
11 Signal Gen~
195 329 388 0 64 64
0 32 31 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1112014848 1133903872 1133903872
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 270
20
1 50 300 300 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
6 0/600V
-22 -30 20 -22
2 V2
-7 -40 7 -32
0
0
40 %D %1 %2 DC 0 SIN(300 300 50 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
1 V
8277 0 0
2
43274.8 0
0
7 Ground~
168 572 305 0 1 3
0 2
0
0 0 53360 180
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3457 0 0
2
43274.7 5
0
2 +V
167 619 325 0 1 3
0 34
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3796 0 0
2
43274.7 4
0
7 Ground~
168 619 401 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6904 0 0
2
43274.7 3
0
10 Op-Amp5:A~
219 619 377 0 5 11
0 28 27 34 2 33
0
0 0 848 0
5 LM358
15 -25 50 -17
2 U1
26 -35 40 -27
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
0
11

0 3 2 7 4 6 3 2 7 4
6 0
88 0 0 0 0 0 0 0
1 U
8602 0 0
2
43274.7 2
0
11 Resistor:A~
219 862 391 0 2 5
0 11 16
0
0 0 880 90
3 56k
8 0 29 8
3 R13
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3607 0 0
2
43274.8 0
0
11 Resistor:A~
219 850 583 0 2 5
0 3 8
0
0 0 880 90
3 56k
8 0 29 8
3 R28
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9456 0 0
2
43274.8 6
0
11 Resistor:A~
219 1010 632 0 2 5
0 5 4
0
0 0 880 180
4 200k
-14 -14 14 -6
3 R27
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3348 0 0
2
43274.8 5
0
11 Resistor:A~
219 964 528 0 3 5
0 2 6 -1
0
0 0 880 270
4 200k
9 1 37 9
3 R10
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7418 0 0
2
43274.8 4
0
11 Resistor:A~
219 905 558 0 2 5
0 8 6
0
0 0 880 0
4 10k2
-14 -14 14 -6
2 R9
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3281 0 0
2
43274.8 3
0
11 Resistor:A~
219 903 605 0 2 5
0 3 4
0
0 0 880 0
4 10k2
-14 -14 14 -6
2 R8
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3613 0 0
2
43274.8 2
0
11 Resistor:A~
219 812 605 0 2 5
0 9 3
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R7
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9506 0 0
2
43274.8 1
0
11 Resistor:A~
219 813 558 0 2 5
0 10 8
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R6
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6773 0 0
2
43274.8 0
0
11 Resistor:A~
219 825 368 0 2 5
0 18 16
0
0 0 880 0
4 224k
-14 -14 14 -6
3 R11
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
8799 0 0
2
43274.8 11
0
11 Resistor:A~
219 824 415 0 2 5
0 17 11
0
0 0 880 0
4 224k
-14 -14 14 -6
3 R12
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7433 0 0
2
43274.8 10
0
11 Resistor:A~
219 915 415 0 2 5
0 11 12
0
0 0 880 0
4 10k2
-13 -14 15 -6
3 R25
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6183 0 0
2
43274.8 9
0
11 Resistor:A~
219 917 368 0 2 5
0 16 14
0
0 0 880 0
4 10k2
-13 -14 15 -6
3 R26
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5243 0 0
2
43274.8 8
0
11 Resistor:A~
219 976 338 0 3 5
0 2 14 -1
0
0 0 880 270
4 200k
9 1 37 9
3 R14
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3217 0 0
2
43274.8 7
0
11 Resistor:A~
219 1022 442 0 2 5
0 13 12
0
0 0 880 180
4 200k
-14 -14 14 -6
3 R15
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
998 0 0
2
43274.8 6
0
11 Resistor:A~
219 570 529 0 3 5
0 2 20 -1
0
0 0 880 270
3 11k
10 1 31 9
3 R24
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9272 0 0
2
43274.8 12
0
11 Resistor:A~
219 616 633 0 2 5
0 25 19
0
0 0 880 180
3 11k
-13 -14 8 -6
3 R23
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3327 0 0
2
43274.8 11
0
11 Resistor:A~
219 441 577 0 2 5
0 22 21
0
0 0 880 90
3 56k
8 0 29 8
3 R22
5 -10 26 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
466 0 0
2
43274.8 10
0
11 Resistor:A~
219 403 600 0 2 5
0 23 22
0
0 0 880 0
4 224k
-14 -14 14 -6
3 R21
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
6854 0 0
2
43274.8 9
0
11 Resistor:A~
219 404 553 0 2 5
0 24 21
0
0 0 880 0
4 224k
-14 -14 14 -6
3 R20
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7745 0 0
2
43274.8 8
0
11 Resistor:A~
219 487 555 0 2 5
0 21 20
0
0 0 880 0
4 124k
-14 -14 14 -6
3 R19
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5764 0 0
2
43274.8 7
0
11 Resistor:A~
219 484 598 0 2 5
0 22 19
0
0 0 880 0
4 124k
-14 -14 14 -6
3 R18
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
5379 0 0
2
43274.8 6
0
11 Resistor:A~
219 486 409 0 2 5
0 30 27
0
0 0 880 0
4 124k
-14 -14 14 -6
3 R17
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7186 0 0
2
43274.8 0
0
11 Resistor:A~
219 489 366 0 2 5
0 29 28
0
0 0 880 0
4 124k
-14 -14 14 -6
3 R16
-10 -24 11 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9136 0 0
2
43274.8 0
0
11 Resistor:A~
219 406 364 0 2 5
0 32 29
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
7143 0 0
2
43274.8 3
0
11 Resistor:A~
219 405 411 0 2 5
0 31 30
0
0 0 880 0
4 224k
-14 -14 14 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9634 0 0
2
43274.8 2
0
11 Resistor:A~
219 443 388 0 2 5
0 30 29
0
0 0 880 90
3 56k
8 0 29 8
2 R5
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
3661 0 0
2
43274.8 1
0
11 Resistor:A~
219 618 444 0 2 5
0 33 27
0
0 0 880 180
4 6.8k
-16 -14 12 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
4323 0 0
2
43274.7 1
0
11 Resistor:A~
219 572 340 0 3 5
0 2 28 -1
0
0 0 880 270
4 6.8k
7 1 35 9
2 R3
8 -10 22 -2
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 0 0 0 0
1 R
9804 0 0
2
43274.7 0
0
56
1 0 3 0 0 4224 0 28 0 0 12 2
885 605
849 605
2 0 4 0 0 4096 0 28 0 0 4 2
921 605
964 605
5 1 5 0 0 8320 0 5 25 0 0 4
1029 564
1044 564
1044 632
1028 632
2 2 4 0 0 8320 0 25 5 0 0 4
992 632
964 632
964 570
993 570
1 1 2 0 0 4224 0 2 26 0 0 2
964 501
964 510
2 0 6 0 0 4224 0 27 0 0 7 2
923 558
964 558
1 2 6 0 0 0 0 5 26 0 0 5
993 558
964 558
964 559
964 559
964 546
1 3 7 0 0 4224 0 3 5 0 0 2
1011 532
1011 551
1 4 2 0 0 0 0 4 5 0 0 2
1011 583
1011 577
1 0 8 0 0 4224 0 27 0 0 11 2
887 558
850 558
2 2 8 0 0 0 0 30 24 0 0 3
831 558
850 558
850 565
2 1 3 0 0 0 0 29 24 0 0 3
830 605
850 605
850 601
1 2 9 0 0 8320 0 29 1 0 0 4
794 605
779 605
779 587
764 587
1 1 10 0 0 8320 0 1 30 0 0 4
764 577
779 577
779 558
795 558
1 0 11 0 0 4224 0 33 0 0 26 2
897 415
861 415
2 0 12 0 0 4096 0 33 0 0 18 2
933 415
976 415
5 1 13 0 0 8320 0 6 36 0 0 4
1041 374
1056 374
1056 442
1040 442
2 2 12 0 0 8320 0 36 6 0 0 4
1004 442
976 442
976 380
1005 380
1 1 2 0 0 0 0 9 35 0 0 2
976 311
976 320
2 0 14 0 0 4224 0 34 0 0 21 2
935 368
976 368
1 2 14 0 0 0 0 6 35 0 0 5
1005 368
976 368
976 369
976 369
976 356
1 3 15 0 0 4224 0 8 6 0 0 2
1023 342
1023 361
1 4 2 0 0 0 0 7 6 0 0 2
1023 393
1023 387
1 0 16 0 0 4224 0 34 0 0 25 2
899 368
862 368
2 2 16 0 0 0 0 31 23 0 0 3
843 368
862 368
862 373
2 1 11 0 0 0 0 32 23 0 0 3
842 415
862 415
862 409
1 2 17 0 0 8320 0 32 10 0 0 4
806 415
791 415
791 397
776 397
1 1 18 0 0 8320 0 10 31 0 0 4
776 387
791 387
791 368
807 368
2 0 19 0 0 4224 0 43 0 0 38 2
502 598
570 598
2 0 20 0 0 4224 0 42 0 0 40 2
505 555
570 555
1 0 21 0 0 8320 0 42 0 0 33 3
469 555
469 553
441 553
1 0 22 0 0 8320 0 43 0 0 34 3
466 598
466 600
441 600
2 2 21 0 0 0 0 41 39 0 0 3
422 553
441 553
441 559
2 1 22 0 0 0 0 40 39 0 0 3
421 600
441 600
441 595
1 2 23 0 0 8320 0 40 15 0 0 4
385 600
370 600
370 582
358 582
1 1 24 0 0 8320 0 15 41 0 0 4
358 572
370 572
370 553
386 553
5 1 25 0 0 8320 0 11 38 0 0 4
635 566
650 566
650 633
634 633
2 2 19 0 0 0 0 38 11 0 0 4
598 633
570 633
570 572
599 572
1 1 2 0 0 128 0 14 37 0 0 2
570 502
570 511
1 2 20 0 0 0 0 11 37 0 0 3
599 560
570 560
570 547
1 3 26 0 0 4224 0 13 11 0 0 2
617 523
617 553
1 4 2 0 0 0 0 12 11 0 0 2
617 584
617 579
2 0 27 0 0 4224 0 44 0 0 52 2
504 409
572 409
2 0 28 0 0 4224 0 45 0 0 54 2
507 366
572 366
1 0 29 0 0 8320 0 45 0 0 47 3
471 366
471 364
443 364
1 0 30 0 0 8320 0 44 0 0 48 3
468 409
468 411
443 411
2 2 29 0 0 0 0 46 48 0 0 3
424 364
443 364
443 370
2 1 30 0 0 0 0 47 48 0 0 3
423 411
443 411
443 406
1 2 31 0 0 8320 0 47 18 0 0 4
387 411
372 411
372 393
360 393
1 1 32 0 0 8320 0 18 46 0 0 4
360 383
372 383
372 364
388 364
5 1 33 0 0 8320 0 22 49 0 0 4
637 377
652 377
652 444
636 444
2 2 27 0 0 128 0 49 22 0 0 4
600 444
572 444
572 383
601 383
1 1 2 0 0 128 0 19 50 0 0 2
572 313
572 322
1 2 28 0 0 0 0 22 50 0 0 3
601 371
572 371
572 358
1 3 34 0 0 4224 0 20 22 0 0 2
619 334
619 364
1 4 2 0 0 0 0 21 22 0 0 2
619 395
619 390
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.1 0.0004 0.0004
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
