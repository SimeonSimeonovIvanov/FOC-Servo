CircuitMaker Text
5.6
Probes: 1
U1A_1
Transient Analysis
0 586 86 65280
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 160 10
176 79 1918 1019
7 5.000 V
7 5.000 V
3 GND
0 0
3 100 0 2 1
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.604255 0.500000
344 175 2086 742
9961490 0
0
6 Title:
5 Name:
0
0
0
19
7 Ground~
168 439 146 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3641 0 0
2
43307 5
0
11 Signal Gen~
195 394 97 0 64 64
0 4 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 1070805811 1068289229
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 266
20
1 1000 1.65 1.35 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
7 300m/3V
-24 -30 25 -22
2 V3
-7 -40 7 -32
0
0
42 %D %1 %2 DC 0 SIN(1.65 1.35 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3104 0 0
2
43307 4
0
2 +V
167 495 106 0 1 3
0 5
0
0 0 53616 90
5 1.65V
-38 -5 -3 3
2 V2
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3296 0 0
2
43307 3
0
7 Ground~
168 534 124 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8534 0 0
2
43307 2
0
2 +V
167 534 70 0 1 3
0 3
0
0 0 53616 0
4 3.3V
-12 -16 16 -8
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
949 0 0
2
43307 1
0
8 Op-Amp5~
219 534 98 0 5 11
0 5 7 3 2 6
0
0 0 848 0
10 LM6132A/NS
8 6 78 14
3 U1A
9 -14 30 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 3 2 8 4 1 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 1 1 0
1 U
3371 0 0
2
43307 0
0
8 Op-Amp5~
219 236 91 0 5 11
0 10 14 12 2 13
0
0 0 848 0
10 LM6132A/NS
8 6 78 14
3 U1B
9 -14 30 -6
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
5 SMD8A
16

0 5 6 8 4 7 3 2 8 4
1 5 6 8 4 7 0
88 0 0 256 2 2 1 0
1 U
7311 0 0
2
43307 6
0
2 +V
167 236 63 0 1 3
0 12
0
0 0 53616 0
4 3.3V
-12 -16 16 -8
2 V4
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3409 0 0
2
43307 5
0
7 Ground~
168 236 117 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3526 0 0
2
43307 4
0
2 +V
167 142 87 0 1 3
0 11
0
0 0 53616 90
5 1.65V
-38 -5 -3 3
2 V5
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4129 0 0
2
43307 3
0
2 +V
167 141 141 0 1 3
0 9
0
0 0 53616 90
4 3.3V
-35 -5 -7 3
2 V7
-7 -25 7 -17
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
6278 0 0
2
43307 2
0
11 Signal Gen~
195 44 102 0 64 64
0 8 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 1065353216 1148846080 0 1068289229
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 18
20
1 1000 0 1.35 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 848 0
11 -1.35/1.35V
-38 -30 39 -22
2 V6
-7 -40 7 -32
0
0
39 %D %1 %2 DC 0 SIN(0 1.35 1k 0 0) AC 1 0
0
0
4 SIP2
5

0 1 2 1 2 0
86 0 0 0 1 0 0 0
1 V
3482 0 0
2
43307 1
0
7 Ground~
168 89 149 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8323 0 0
2
43307 0
0
11 Resistor:A~
219 534 35 0 2 5
0 7 6
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R2
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3984 0 0
2
43307 7
0
11 Resistor:A~
219 478 92 0 2 5
0 4 7
0
0 0 880 0
2 5k
-7 -14 7 -6
2 R1
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7622 0 0
2
43307 6
0
11 Resistor:A~
219 180 85 0 3 5
0 11 14 1
0
0 0 880 0
4 3.3k
-14 -14 14 -6
2 R3
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
816 0 0
2
43307 10
0
11 Resistor:A~
219 236 28 0 2 5
0 14 13
0
0 0 880 0
4 3.3k
-14 -14 14 -6
2 R4
-7 -24 7 -16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
4656 0 0
2
43307 9
0
11 Resistor:A~
219 180 97 0 2 5
0 8 10
0
0 0 880 0
4 3.3k
-13 19 15 27
2 R5
-12 8 2 16
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
6356 0 0
2
43307 8
0
11 Resistor:A~
219 180 139 0 4 5
0 10 9 0 1
0
0 0 880 180
4 3.3k
-14 18 14 26
2 R6
-11 7 3 15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
7479 0 0
2
43307 7
0
19
1 3 3 0 0 4240 0 5 6 0 0 2
534 79
534 85
1 2 2 0 0 4240 0 1 2 0 0 3
439 140
439 102
425 102
1 1 4 0 0 4240 0 2 15 0 0 2
425 92
460 92
1 1 5 0 0 4240 0 3 6 0 0 2
506 104
516 104
1 4 2 0 0 16 0 4 6 0 0 2
534 118
534 111
2 5 6 0 0 8336 0 14 6 0 0 4
552 35
585 35
585 98
552 98
1 0 7 0 0 8336 0 14 0 0 8 3
516 35
504 35
504 92
2 2 7 0 0 16 0 15 6 0 0 2
496 92
516 92
1 1 8 0 0 4224 0 18 12 0 0 2
162 97
75 97
1 2 2 0 0 0 0 13 12 0 0 3
89 143
89 107
75 107
1 2 9 0 0 4224 0 11 19 0 0 2
152 139
162 139
1 0 10 0 0 8320 0 19 0 0 13 3
198 139
206 139
206 97
2 1 10 0 0 0 0 18 7 0 0 2
198 97
218 97
1 1 11 0 0 4224 0 10 16 0 0 2
153 85
162 85
1 3 12 0 0 4224 0 8 7 0 0 2
236 72
236 78
1 4 2 0 0 0 0 9 7 0 0 2
236 111
236 104
2 5 13 0 0 8320 0 17 7 0 0 4
254 28
287 28
287 91
254 91
1 0 14 0 0 8320 0 17 0 0 19 3
218 28
206 28
206 85
2 2 14 0 0 0 0 16 7 0 0 2
198 85
218 85
0
0
2065 0 1
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0.005 2e-05 2e-05
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
